module testbench_scaled;

    //neuron addresses
        source_addresses[129] = 12'd1153;        source_addresses[155] = 12'd1179;        source_addresses[156] = 12'd1180;        source_addresses[157] = 12'd1181;        source_addresses[158] = 12'd1182;        source_addresses[159] = 12'd1183;        source_addresses[182] = 12'd1206;        source_addresses[183] = 12'd1207;        source_addresses[184] = 12'd1208;        source_addresses[185] = 12'd1209;        source_addresses[186] = 12'd1210;        source_addresses[187] = 12'd1211;        source_addresses[209] = 12'd1233;        source_addresses[210] = 12'd1234;        source_addresses[211] = 12'd1235;        source_addresses[212] = 12'd1236;        source_addresses[213] = 12'd1237;        source_addresses[215] = 12'd1239;        source_addresses[216] = 12'd1240;        source_addresses[236] = 12'd1260;        source_addresses[237] = 12'd1261;        source_addresses[238] = 12'd1262;        source_addresses[239] = 12'd1263;        source_addresses[240] = 12'd1264;        source_addresses[241] = 12'd1265;        source_addresses[244] = 12'd1268;        source_addresses[263] = 12'd1287;        source_addresses[264] = 12'd1288;        source_addresses[265] = 12'd1289;        source_addresses[268] = 12'd1292;        source_addresses[269] = 12'd1293;        source_addresses[272] = 12'd1296;        source_addresses[290] = 12'd1314;        source_addresses[291] = 12'd1315;        source_addresses[292] = 12'd1316;        source_addresses[300] = 12'd1324;
        source_addresses[301] = 12'd1325;        source_addresses[318] = 12'd1342;        source_addresses[319] = 12'd1343;        source_addresses[320] = 12'd1344;        source_addresses[328] = 12'd1352;        source_addresses[329] = 12'd1353;        source_addresses[345] = 12'd1369;        source_addresses[346] = 12'd1370;        source_addresses[356] = 12'd1380;        source_addresses[357] = 12'd1381;        source_addresses[358] = 12'd1382;        source_addresses[372] = 12'd1396;        source_addresses[373] = 12'd1397;        source_addresses[384] = 12'd1408;        source_addresses[385] = 12'd1409;        source_addresses[386] = 12'd1410;        source_addresses[399] = 12'd1423;        source_addresses[400] = 12'd1424;
        source_addresses[412] = 12'd1436;        source_addresses[413] = 12'd1437;        source_addresses[414] = 12'd1438;        source_addresses[427] = 12'd1451;        source_addresses[428] = 12'd1452;        source_addresses[440] = 12'd1464;        source_addresses[441] = 12'd1465;        source_addresses[455] = 12'd1479;        source_addresses[456] = 12'd1480;        source_addresses[468] = 12'd1492;        source_addresses[483] = 12'd1507;        source_addresses[484] = 12'd1508;        source_addresses[495] = 12'd1519;        source_addresses[496] = 12'd1520;        source_addresses[511] = 12'd1535;        source_addresses[522] = 12'd1546;        source_addresses[539] = 12'd1563;        source_addresses[540] = 12'd1564;        source_addresses[548] = 12'd1572;        source_addresses[549] = 12'd1573;        source_addresses[567] = 12'd1591;        source_addresses[568] = 12'd1592;        source_addresses[574] = 12'd1598;        source_addresses[575] = 12'd1599;        source_addresses[576] = 12'd1600;        source_addresses[595] = 12'd1619;        source_addresses[596] = 12'd1620;        source_addresses[597] = 12'd1621;        source_addresses[598] = 12'd1622;        source_addresses[599] = 12'd1623;        source_addresses[600] = 12'd1624;
        source_addresses[601] = 12'd1625;        source_addresses[602] = 12'd1626;        source_addresses[603] = 12'd1627;        source_addresses[623] = 12'd1647;        source_addresses[624] = 12'd1648;        source_addresses[625] = 12'd1649;        source_addresses[626] = 12'd1650;        source_addresses[627] = 12'd1651;        source_addresses[628] = 12'd1652;        source_addresses[629] = 12'd1653;        source_addresses[653] = 12'd1677;        source_addresses[654] = 12'd1678;        source_addresses[655] = 12'd1679;