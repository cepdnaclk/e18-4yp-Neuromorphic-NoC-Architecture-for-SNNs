module adder(
    input wire [31:0] weight, 
    input wire [31:0] decayed_potential, 
    output reg [31:0] potential, 
    output reg spike);

    // Addition and comparison
    
     



endmodule