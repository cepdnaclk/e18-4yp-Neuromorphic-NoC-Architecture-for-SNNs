// MAC unit can process 4 input spikes together
// 4 spike inputs  
// 4 weights corresponding to the synapse

/*  Floating point addition
    Moving through the next four connections ?*/
`timescale 1ns/100ps
// `include "Addition_Subtraction.v"


module mac(
    
    input wire CLK,                             //input clock
    input wire[11:0] neuron_address,            //neuron address
    input wire[11:0] source_address,            //source address of 12 bits
    input wire[weights_array_width-1:0] weights_array,            //weights array used during intialization 32x5=160 bits
    input wire[number_of_connections*number_of_address_bits-1:0] source_addresses_array,          //corresponding source address array used during initialization 12x5=60 bits
    input wire clear,                       //signal to signify the end of the timestep
    output reg[31:0] mult_output               //output of 32 bits to the adder
    );             

    parameter number_of_connections = 784;
    parameter number_of_address_bits = 12;
    parameter number_of_units = 1024;
    parameter weights_array_width = 32 * number_of_connections;

    integer i;                      //iterate through for the sources addresses
    integer index;                  //get array index of the connection
    reg incoming_spikes[0:number_of_connections-1];   //note incoming spikes
    reg spikes[0:number_of_connections-1];            //received stored spikes
    reg[31:0] weights [0:number_of_connections-1];    //array to store 5 weights
    reg[11:0] source_addresses [0:number_of_connections-1];    //array to store corresponding 5 source addresses
    reg break;
    reg[31:0] accumulated_weight;   //get the accumulated weight
    reg[31:0] considered_weight;    //weight to be added
    wire[31:0] added_weight;         //weight
    wire exception;                 //addition exception
    integer topBorder;
    integer lowerBorder;

    //addition block to add weights
    Addition_Subtraction add1(accumulated_weight, considered_weight, 1'b0, excpetion, added_weight);

    always @(weights_array, source_addresses_array) begin
        //break up the weights
        weights[0]=weights_array[25087:25056];      weights[1]=weights_array[25055:25024];      weights[2]=weights_array[25023:24992];      weights[3]=weights_array[24991:24960];      weights[4]=weights_array[24959:24928];      weights[5]=weights_array[24927:24896];      weights[6]=weights_array[24895:24864];      weights[7]=weights_array[24863:24832];      weights[8]=weights_array[24831:24800];      weights[9]=weights_array[24799:24768];      weights[10]=weights_array[24767:24736];      weights[11]=weights_array[24735:24704];      weights[12]=weights_array[24703:24672];      weights[13]=weights_array[24671:24640];      weights[14]=weights_array[24639:24608];      weights[15]=weights_array[24607:24576];      weights[16]=weights_array[24575:24544];      weights[17]=weights_array[24543:24512];      weights[18]=weights_array[24511:24480];      weights[19]=weights_array[24479:24448];      weights[20]=weights_array[24447:24416];      weights[21]=weights_array[24415:24384];      weights[22]=weights_array[24383:24352];      weights[23]=weights_array[24351:24320];      weights[24]=weights_array[24319:24288];      weights[25]=weights_array[24287:24256];      weights[26]=weights_array[24255:24224];      weights[27]=weights_array[24223:24192];      weights[28]=weights_array[24191:24160];      weights[29]=weights_array[24159:24128];      weights[30]=weights_array[24127:24096];      weights[31]=weights_array[24095:24064];      weights[32]=weights_array[24063:24032];      weights[33]=weights_array[24031:24000];      weights[34]=weights_array[23999:23968];      weights[35]=weights_array[23967:23936];      weights[36]=weights_array[23935:23904];      weights[37]=weights_array[23903:23872];      weights[38]=weights_array[23871:23840];      weights[39]=weights_array[23839:23808];      weights[40]=weights_array[23807:23776];      weights[41]=weights_array[23775:23744];      weights[42]=weights_array[23743:23712];      weights[43]=weights_array[23711:23680];      weights[44]=weights_array[23679:23648];      weights[45]=weights_array[23647:23616];      weights[46]=weights_array[23615:23584];      weights[47]=weights_array[23583:23552];      weights[48]=weights_array[23551:23520];      weights[49]=weights_array[23519:23488];      weights[50]=weights_array[23487:23456];      weights[51]=weights_array[23455:23424];      weights[52]=weights_array[23423:23392];      weights[53]=weights_array[23391:23360];      weights[54]=weights_array[23359:23328];      weights[55]=weights_array[23327:23296];      weights[56]=weights_array[23295:23264];      weights[57]=weights_array[23263:23232];      weights[58]=weights_array[23231:23200];      weights[59]=weights_array[23199:23168];      weights[60]=weights_array[23167:23136];      weights[61]=weights_array[23135:23104];      weights[62]=weights_array[23103:23072];      weights[63]=weights_array[23071:23040];      weights[64]=weights_array[23039:23008];      weights[65]=weights_array[23007:22976];      weights[66]=weights_array[22975:22944];      weights[67]=weights_array[22943:22912];      weights[68]=weights_array[22911:22880];      weights[69]=weights_array[22879:22848];      weights[70]=weights_array[22847:22816];      weights[71]=weights_array[22815:22784];      weights[72]=weights_array[22783:22752];      weights[73]=weights_array[22751:22720];      weights[74]=weights_array[22719:22688];      weights[75]=weights_array[22687:22656];      weights[76]=weights_array[22655:22624];      weights[77]=weights_array[22623:22592];      weights[78]=weights_array[22591:22560];      weights[79]=weights_array[22559:22528];      weights[80]=weights_array[22527:22496];      weights[81]=weights_array[22495:22464];      weights[82]=weights_array[22463:22432];      weights[83]=weights_array[22431:22400];      weights[84]=weights_array[22399:22368];      weights[85]=weights_array[22367:22336];      weights[86]=weights_array[22335:22304];      weights[87]=weights_array[22303:22272];      weights[88]=weights_array[22271:22240];      weights[89]=weights_array[22239:22208];      weights[90]=weights_array[22207:22176];      weights[91]=weights_array[22175:22144];      weights[92]=weights_array[22143:22112];      weights[93]=weights_array[22111:22080];      weights[94]=weights_array[22079:22048];      weights[95]=weights_array[22047:22016];      weights[96]=weights_array[22015:21984];      weights[97]=weights_array[21983:21952];      weights[98]=weights_array[21951:21920];      weights[99]=weights_array[21919:21888];      weights[100]=weights_array[21887:21856];      weights[101]=weights_array[21855:21824];      weights[102]=weights_array[21823:21792];      weights[103]=weights_array[21791:21760];      weights[104]=weights_array[21759:21728];      weights[105]=weights_array[21727:21696];      weights[106]=weights_array[21695:21664];      weights[107]=weights_array[21663:21632];      weights[108]=weights_array[21631:21600];      weights[109]=weights_array[21599:21568];      weights[110]=weights_array[21567:21536];      weights[111]=weights_array[21535:21504];      weights[112]=weights_array[21503:21472];      weights[113]=weights_array[21471:21440];      weights[114]=weights_array[21439:21408];      weights[115]=weights_array[21407:21376];      weights[116]=weights_array[21375:21344];      weights[117]=weights_array[21343:21312];      weights[118]=weights_array[21311:21280];      weights[119]=weights_array[21279:21248];      weights[120]=weights_array[21247:21216];      weights[121]=weights_array[21215:21184];      weights[122]=weights_array[21183:21152];      weights[123]=weights_array[21151:21120];      weights[124]=weights_array[21119:21088];      weights[125]=weights_array[21087:21056];      weights[126]=weights_array[21055:21024];      weights[127]=weights_array[21023:20992];      weights[128]=weights_array[20991:20960];      weights[129]=weights_array[20959:20928];      weights[130]=weights_array[20927:20896];      weights[131]=weights_array[20895:20864];      weights[132]=weights_array[20863:20832];      weights[133]=weights_array[20831:20800];      weights[134]=weights_array[20799:20768];      weights[135]=weights_array[20767:20736];      weights[136]=weights_array[20735:20704];      weights[137]=weights_array[20703:20672];      weights[138]=weights_array[20671:20640];      weights[139]=weights_array[20639:20608];      weights[140]=weights_array[20607:20576];      weights[141]=weights_array[20575:20544];      weights[142]=weights_array[20543:20512];      weights[143]=weights_array[20511:20480];      weights[144]=weights_array[20479:20448];      weights[145]=weights_array[20447:20416];      weights[146]=weights_array[20415:20384];      weights[147]=weights_array[20383:20352];      weights[148]=weights_array[20351:20320];      weights[149]=weights_array[20319:20288];      weights[150]=weights_array[20287:20256];      weights[151]=weights_array[20255:20224];      weights[152]=weights_array[20223:20192];      weights[153]=weights_array[20191:20160];      weights[154]=weights_array[20159:20128];      weights[155]=weights_array[20127:20096];      weights[156]=weights_array[20095:20064];      weights[157]=weights_array[20063:20032];      weights[158]=weights_array[20031:20000];      weights[159]=weights_array[19999:19968];      weights[160]=weights_array[19967:19936];      weights[161]=weights_array[19935:19904];      weights[162]=weights_array[19903:19872];      weights[163]=weights_array[19871:19840];      weights[164]=weights_array[19839:19808];      weights[165]=weights_array[19807:19776];      weights[166]=weights_array[19775:19744];      weights[167]=weights_array[19743:19712];      weights[168]=weights_array[19711:19680];      weights[169]=weights_array[19679:19648];      weights[170]=weights_array[19647:19616];      weights[171]=weights_array[19615:19584];      weights[172]=weights_array[19583:19552];      weights[173]=weights_array[19551:19520];      weights[174]=weights_array[19519:19488];      weights[175]=weights_array[19487:19456];      weights[176]=weights_array[19455:19424];      weights[177]=weights_array[19423:19392];      weights[178]=weights_array[19391:19360];      weights[179]=weights_array[19359:19328];      weights[180]=weights_array[19327:19296];      weights[181]=weights_array[19295:19264];      weights[182]=weights_array[19263:19232];      weights[183]=weights_array[19231:19200];      weights[184]=weights_array[19199:19168];      weights[185]=weights_array[19167:19136];      weights[186]=weights_array[19135:19104];      weights[187]=weights_array[19103:19072];      weights[188]=weights_array[19071:19040];      weights[189]=weights_array[19039:19008];      weights[190]=weights_array[19007:18976];      weights[191]=weights_array[18975:18944];      weights[192]=weights_array[18943:18912];      weights[193]=weights_array[18911:18880];      weights[194]=weights_array[18879:18848];      weights[195]=weights_array[18847:18816];      weights[196]=weights_array[18815:18784];      weights[197]=weights_array[18783:18752];      weights[198]=weights_array[18751:18720];      weights[199]=weights_array[18719:18688];      weights[200]=weights_array[18687:18656];      weights[201]=weights_array[18655:18624];      weights[202]=weights_array[18623:18592];      weights[203]=weights_array[18591:18560];      weights[204]=weights_array[18559:18528];      weights[205]=weights_array[18527:18496];      weights[206]=weights_array[18495:18464];      weights[207]=weights_array[18463:18432];      weights[208]=weights_array[18431:18400];      weights[209]=weights_array[18399:18368];      weights[210]=weights_array[18367:18336];      weights[211]=weights_array[18335:18304];      weights[212]=weights_array[18303:18272];      weights[213]=weights_array[18271:18240];      weights[214]=weights_array[18239:18208];      weights[215]=weights_array[18207:18176];      weights[216]=weights_array[18175:18144];      weights[217]=weights_array[18143:18112];      weights[218]=weights_array[18111:18080];      weights[219]=weights_array[18079:18048];      weights[220]=weights_array[18047:18016];      weights[221]=weights_array[18015:17984];      weights[222]=weights_array[17983:17952];      weights[223]=weights_array[17951:17920];      weights[224]=weights_array[17919:17888];      weights[225]=weights_array[17887:17856];      weights[226]=weights_array[17855:17824];      weights[227]=weights_array[17823:17792];      weights[228]=weights_array[17791:17760];      weights[229]=weights_array[17759:17728];      weights[230]=weights_array[17727:17696];      weights[231]=weights_array[17695:17664];      weights[232]=weights_array[17663:17632];      weights[233]=weights_array[17631:17600];      weights[234]=weights_array[17599:17568];      weights[235]=weights_array[17567:17536];      weights[236]=weights_array[17535:17504];      weights[237]=weights_array[17503:17472];      weights[238]=weights_array[17471:17440];      weights[239]=weights_array[17439:17408];      weights[240]=weights_array[17407:17376];      weights[241]=weights_array[17375:17344];      weights[242]=weights_array[17343:17312];      weights[243]=weights_array[17311:17280];      weights[244]=weights_array[17279:17248];      weights[245]=weights_array[17247:17216];      weights[246]=weights_array[17215:17184];      weights[247]=weights_array[17183:17152];      weights[248]=weights_array[17151:17120];      weights[249]=weights_array[17119:17088];      weights[250]=weights_array[17087:17056];      weights[251]=weights_array[17055:17024];      weights[252]=weights_array[17023:16992];      weights[253]=weights_array[16991:16960];      weights[254]=weights_array[16959:16928];      weights[255]=weights_array[16927:16896];      weights[256]=weights_array[16895:16864];      weights[257]=weights_array[16863:16832];      weights[258]=weights_array[16831:16800];      weights[259]=weights_array[16799:16768];      weights[260]=weights_array[16767:16736];      weights[261]=weights_array[16735:16704];      weights[262]=weights_array[16703:16672];      weights[263]=weights_array[16671:16640];      weights[264]=weights_array[16639:16608];      weights[265]=weights_array[16607:16576];      weights[266]=weights_array[16575:16544];      weights[267]=weights_array[16543:16512];      weights[268]=weights_array[16511:16480];      weights[269]=weights_array[16479:16448];      weights[270]=weights_array[16447:16416];      weights[271]=weights_array[16415:16384];      weights[272]=weights_array[16383:16352];      weights[273]=weights_array[16351:16320];      weights[274]=weights_array[16319:16288];      weights[275]=weights_array[16287:16256];      weights[276]=weights_array[16255:16224];      weights[277]=weights_array[16223:16192];      weights[278]=weights_array[16191:16160];      weights[279]=weights_array[16159:16128];      weights[280]=weights_array[16127:16096];      weights[281]=weights_array[16095:16064];      weights[282]=weights_array[16063:16032];      weights[283]=weights_array[16031:16000];      weights[284]=weights_array[15999:15968];      weights[285]=weights_array[15967:15936];      weights[286]=weights_array[15935:15904];      weights[287]=weights_array[15903:15872];      weights[288]=weights_array[15871:15840];      weights[289]=weights_array[15839:15808];      weights[290]=weights_array[15807:15776];      weights[291]=weights_array[15775:15744];      weights[292]=weights_array[15743:15712];      weights[293]=weights_array[15711:15680];      weights[294]=weights_array[15679:15648];      weights[295]=weights_array[15647:15616];      weights[296]=weights_array[15615:15584];      weights[297]=weights_array[15583:15552];      weights[298]=weights_array[15551:15520];      weights[299]=weights_array[15519:15488];      weights[300]=weights_array[15487:15456];      weights[301]=weights_array[15455:15424];      weights[302]=weights_array[15423:15392];      weights[303]=weights_array[15391:15360];      weights[304]=weights_array[15359:15328];      weights[305]=weights_array[15327:15296];      weights[306]=weights_array[15295:15264];      weights[307]=weights_array[15263:15232];      weights[308]=weights_array[15231:15200];      weights[309]=weights_array[15199:15168];      weights[310]=weights_array[15167:15136];      weights[311]=weights_array[15135:15104];      weights[312]=weights_array[15103:15072];      weights[313]=weights_array[15071:15040];      weights[314]=weights_array[15039:15008];      weights[315]=weights_array[15007:14976];      weights[316]=weights_array[14975:14944];      weights[317]=weights_array[14943:14912];      weights[318]=weights_array[14911:14880];      weights[319]=weights_array[14879:14848];      weights[320]=weights_array[14847:14816];      weights[321]=weights_array[14815:14784];      weights[322]=weights_array[14783:14752];      weights[323]=weights_array[14751:14720];      weights[324]=weights_array[14719:14688];      weights[325]=weights_array[14687:14656];      weights[326]=weights_array[14655:14624];      weights[327]=weights_array[14623:14592];      weights[328]=weights_array[14591:14560];      weights[329]=weights_array[14559:14528];      weights[330]=weights_array[14527:14496];      weights[331]=weights_array[14495:14464];      weights[332]=weights_array[14463:14432];      weights[333]=weights_array[14431:14400];      weights[334]=weights_array[14399:14368];      weights[335]=weights_array[14367:14336];      weights[336]=weights_array[14335:14304];      weights[337]=weights_array[14303:14272];      weights[338]=weights_array[14271:14240];      weights[339]=weights_array[14239:14208];      weights[340]=weights_array[14207:14176];      weights[341]=weights_array[14175:14144];      weights[342]=weights_array[14143:14112];      weights[343]=weights_array[14111:14080];      weights[344]=weights_array[14079:14048];      weights[345]=weights_array[14047:14016];      weights[346]=weights_array[14015:13984];      weights[347]=weights_array[13983:13952];      weights[348]=weights_array[13951:13920];      weights[349]=weights_array[13919:13888];      weights[350]=weights_array[13887:13856];      weights[351]=weights_array[13855:13824];      weights[352]=weights_array[13823:13792];      weights[353]=weights_array[13791:13760];      weights[354]=weights_array[13759:13728];      weights[355]=weights_array[13727:13696];      weights[356]=weights_array[13695:13664];      weights[357]=weights_array[13663:13632];      weights[358]=weights_array[13631:13600];      weights[359]=weights_array[13599:13568];      weights[360]=weights_array[13567:13536];      weights[361]=weights_array[13535:13504];      weights[362]=weights_array[13503:13472];      weights[363]=weights_array[13471:13440];      weights[364]=weights_array[13439:13408];      weights[365]=weights_array[13407:13376];      weights[366]=weights_array[13375:13344];      weights[367]=weights_array[13343:13312];      weights[368]=weights_array[13311:13280];      weights[369]=weights_array[13279:13248];      weights[370]=weights_array[13247:13216];      weights[371]=weights_array[13215:13184];      weights[372]=weights_array[13183:13152];      weights[373]=weights_array[13151:13120];      weights[374]=weights_array[13119:13088];      weights[375]=weights_array[13087:13056];      weights[376]=weights_array[13055:13024];      weights[377]=weights_array[13023:12992];      weights[378]=weights_array[12991:12960];      weights[379]=weights_array[12959:12928];      weights[380]=weights_array[12927:12896];      weights[381]=weights_array[12895:12864];      weights[382]=weights_array[12863:12832];      weights[383]=weights_array[12831:12800];      weights[384]=weights_array[12799:12768];      weights[385]=weights_array[12767:12736];      weights[386]=weights_array[12735:12704];      weights[387]=weights_array[12703:12672];      weights[388]=weights_array[12671:12640];      weights[389]=weights_array[12639:12608];      weights[390]=weights_array[12607:12576];      weights[391]=weights_array[12575:12544];      weights[392]=weights_array[12543:12512];      weights[393]=weights_array[12511:12480];      weights[394]=weights_array[12479:12448];      weights[395]=weights_array[12447:12416];      weights[396]=weights_array[12415:12384];      weights[397]=weights_array[12383:12352];      weights[398]=weights_array[12351:12320];      weights[399]=weights_array[12319:12288];      weights[400]=weights_array[12287:12256];      weights[401]=weights_array[12255:12224];      weights[402]=weights_array[12223:12192];      weights[403]=weights_array[12191:12160];      weights[404]=weights_array[12159:12128];      weights[405]=weights_array[12127:12096];      weights[406]=weights_array[12095:12064];      weights[407]=weights_array[12063:12032];      weights[408]=weights_array[12031:12000];      weights[409]=weights_array[11999:11968];      weights[410]=weights_array[11967:11936];      weights[411]=weights_array[11935:11904];      weights[412]=weights_array[11903:11872];      weights[413]=weights_array[11871:11840];      weights[414]=weights_array[11839:11808];      weights[415]=weights_array[11807:11776];      weights[416]=weights_array[11775:11744];      weights[417]=weights_array[11743:11712];      weights[418]=weights_array[11711:11680];      weights[419]=weights_array[11679:11648];      weights[420]=weights_array[11647:11616];      weights[421]=weights_array[11615:11584];      weights[422]=weights_array[11583:11552];      weights[423]=weights_array[11551:11520];      weights[424]=weights_array[11519:11488];      weights[425]=weights_array[11487:11456];      weights[426]=weights_array[11455:11424];      weights[427]=weights_array[11423:11392];      weights[428]=weights_array[11391:11360];      weights[429]=weights_array[11359:11328];      weights[430]=weights_array[11327:11296];      weights[431]=weights_array[11295:11264];      weights[432]=weights_array[11263:11232];      weights[433]=weights_array[11231:11200];      weights[434]=weights_array[11199:11168];      weights[435]=weights_array[11167:11136];      weights[436]=weights_array[11135:11104];      weights[437]=weights_array[11103:11072];      weights[438]=weights_array[11071:11040];      weights[439]=weights_array[11039:11008];      weights[440]=weights_array[11007:10976];      weights[441]=weights_array[10975:10944];      weights[442]=weights_array[10943:10912];      weights[443]=weights_array[10911:10880];      weights[444]=weights_array[10879:10848];      weights[445]=weights_array[10847:10816];      weights[446]=weights_array[10815:10784];      weights[447]=weights_array[10783:10752];      weights[448]=weights_array[10751:10720];      weights[449]=weights_array[10719:10688];      weights[450]=weights_array[10687:10656];      weights[451]=weights_array[10655:10624];      weights[452]=weights_array[10623:10592];      weights[453]=weights_array[10591:10560];      weights[454]=weights_array[10559:10528];      weights[455]=weights_array[10527:10496];      weights[456]=weights_array[10495:10464];      weights[457]=weights_array[10463:10432];      weights[458]=weights_array[10431:10400];      weights[459]=weights_array[10399:10368];      weights[460]=weights_array[10367:10336];      weights[461]=weights_array[10335:10304];      weights[462]=weights_array[10303:10272];      weights[463]=weights_array[10271:10240];      weights[464]=weights_array[10239:10208];      weights[465]=weights_array[10207:10176];      weights[466]=weights_array[10175:10144];      weights[467]=weights_array[10143:10112];      weights[468]=weights_array[10111:10080];      weights[469]=weights_array[10079:10048];      weights[470]=weights_array[10047:10016];      weights[471]=weights_array[10015:9984];      weights[472]=weights_array[9983:9952];      weights[473]=weights_array[9951:9920];      weights[474]=weights_array[9919:9888];      weights[475]=weights_array[9887:9856];      weights[476]=weights_array[9855:9824];      weights[477]=weights_array[9823:9792];      weights[478]=weights_array[9791:9760];      weights[479]=weights_array[9759:9728];      weights[480]=weights_array[9727:9696];      weights[481]=weights_array[9695:9664];      weights[482]=weights_array[9663:9632];      weights[483]=weights_array[9631:9600];      weights[484]=weights_array[9599:9568];      weights[485]=weights_array[9567:9536];      weights[486]=weights_array[9535:9504];      weights[487]=weights_array[9503:9472];      weights[488]=weights_array[9471:9440];      weights[489]=weights_array[9439:9408];      weights[490]=weights_array[9407:9376];      weights[491]=weights_array[9375:9344];      weights[492]=weights_array[9343:9312];      weights[493]=weights_array[9311:9280];      weights[494]=weights_array[9279:9248];      weights[495]=weights_array[9247:9216];      weights[496]=weights_array[9215:9184];      weights[497]=weights_array[9183:9152];      weights[498]=weights_array[9151:9120];      weights[499]=weights_array[9119:9088];      weights[500]=weights_array[9087:9056];      weights[501]=weights_array[9055:9024];      weights[502]=weights_array[9023:8992];      weights[503]=weights_array[8991:8960];      weights[504]=weights_array[8959:8928];      weights[505]=weights_array[8927:8896];      weights[506]=weights_array[8895:8864];      weights[507]=weights_array[8863:8832];      weights[508]=weights_array[8831:8800];      weights[509]=weights_array[8799:8768];      weights[510]=weights_array[8767:8736];      weights[511]=weights_array[8735:8704];      weights[512]=weights_array[8703:8672];      weights[513]=weights_array[8671:8640];      weights[514]=weights_array[8639:8608];      weights[515]=weights_array[8607:8576];      weights[516]=weights_array[8575:8544];      weights[517]=weights_array[8543:8512];      weights[518]=weights_array[8511:8480];      weights[519]=weights_array[8479:8448];      weights[520]=weights_array[8447:8416];      weights[521]=weights_array[8415:8384];      weights[522]=weights_array[8383:8352];      weights[523]=weights_array[8351:8320];      weights[524]=weights_array[8319:8288];      weights[525]=weights_array[8287:8256];      weights[526]=weights_array[8255:8224];      weights[527]=weights_array[8223:8192];      weights[528]=weights_array[8191:8160];      weights[529]=weights_array[8159:8128];      weights[530]=weights_array[8127:8096];      weights[531]=weights_array[8095:8064];      weights[532]=weights_array[8063:8032];      weights[533]=weights_array[8031:8000];      weights[534]=weights_array[7999:7968];      weights[535]=weights_array[7967:7936];      weights[536]=weights_array[7935:7904];      weights[537]=weights_array[7903:7872];      weights[538]=weights_array[7871:7840];      weights[539]=weights_array[7839:7808];      weights[540]=weights_array[7807:7776];      weights[541]=weights_array[7775:7744];      weights[542]=weights_array[7743:7712];      weights[543]=weights_array[7711:7680];      weights[544]=weights_array[7679:7648];      weights[545]=weights_array[7647:7616];      weights[546]=weights_array[7615:7584];      weights[547]=weights_array[7583:7552];      weights[548]=weights_array[7551:7520];      weights[549]=weights_array[7519:7488];      weights[550]=weights_array[7487:7456];      weights[551]=weights_array[7455:7424];      weights[552]=weights_array[7423:7392];      weights[553]=weights_array[7391:7360];      weights[554]=weights_array[7359:7328];      weights[555]=weights_array[7327:7296];      weights[556]=weights_array[7295:7264];      weights[557]=weights_array[7263:7232];      weights[558]=weights_array[7231:7200];      weights[559]=weights_array[7199:7168];      weights[560]=weights_array[7167:7136];      weights[561]=weights_array[7135:7104];      weights[562]=weights_array[7103:7072];      weights[563]=weights_array[7071:7040];      weights[564]=weights_array[7039:7008];      weights[565]=weights_array[7007:6976];      weights[566]=weights_array[6975:6944];      weights[567]=weights_array[6943:6912];      weights[568]=weights_array[6911:6880];      weights[569]=weights_array[6879:6848];      weights[570]=weights_array[6847:6816];      weights[571]=weights_array[6815:6784];      weights[572]=weights_array[6783:6752];      weights[573]=weights_array[6751:6720];      weights[574]=weights_array[6719:6688];      weights[575]=weights_array[6687:6656];      weights[576]=weights_array[6655:6624];      weights[577]=weights_array[6623:6592];      weights[578]=weights_array[6591:6560];      weights[579]=weights_array[6559:6528];      weights[580]=weights_array[6527:6496];      weights[581]=weights_array[6495:6464];      weights[582]=weights_array[6463:6432];      weights[583]=weights_array[6431:6400];      weights[584]=weights_array[6399:6368];      weights[585]=weights_array[6367:6336];      weights[586]=weights_array[6335:6304];      weights[587]=weights_array[6303:6272];      weights[588]=weights_array[6271:6240];      weights[589]=weights_array[6239:6208];      weights[590]=weights_array[6207:6176];      weights[591]=weights_array[6175:6144];      weights[592]=weights_array[6143:6112];      weights[593]=weights_array[6111:6080];      weights[594]=weights_array[6079:6048];      weights[595]=weights_array[6047:6016];      weights[596]=weights_array[6015:5984];      weights[597]=weights_array[5983:5952];      weights[598]=weights_array[5951:5920];      weights[599]=weights_array[5919:5888];      weights[600]=weights_array[5887:5856];      weights[601]=weights_array[5855:5824];      weights[602]=weights_array[5823:5792];      weights[603]=weights_array[5791:5760];      weights[604]=weights_array[5759:5728];      weights[605]=weights_array[5727:5696];      weights[606]=weights_array[5695:5664];      weights[607]=weights_array[5663:5632];      weights[608]=weights_array[5631:5600];      weights[609]=weights_array[5599:5568];      weights[610]=weights_array[5567:5536];      weights[611]=weights_array[5535:5504];      weights[612]=weights_array[5503:5472];      weights[613]=weights_array[5471:5440];      weights[614]=weights_array[5439:5408];      weights[615]=weights_array[5407:5376];      weights[616]=weights_array[5375:5344];      weights[617]=weights_array[5343:5312];      weights[618]=weights_array[5311:5280];      weights[619]=weights_array[5279:5248];      weights[620]=weights_array[5247:5216];      weights[621]=weights_array[5215:5184];      weights[622]=weights_array[5183:5152];      weights[623]=weights_array[5151:5120];      weights[624]=weights_array[5119:5088];      weights[625]=weights_array[5087:5056];      weights[626]=weights_array[5055:5024];      weights[627]=weights_array[5023:4992];      weights[628]=weights_array[4991:4960];      weights[629]=weights_array[4959:4928];      weights[630]=weights_array[4927:4896];      weights[631]=weights_array[4895:4864];      weights[632]=weights_array[4863:4832];      weights[633]=weights_array[4831:4800];      weights[634]=weights_array[4799:4768];      weights[635]=weights_array[4767:4736];      weights[636]=weights_array[4735:4704];      weights[637]=weights_array[4703:4672];      weights[638]=weights_array[4671:4640];      weights[639]=weights_array[4639:4608];      weights[640]=weights_array[4607:4576];      weights[641]=weights_array[4575:4544];      weights[642]=weights_array[4543:4512];      weights[643]=weights_array[4511:4480];      weights[644]=weights_array[4479:4448];      weights[645]=weights_array[4447:4416];      weights[646]=weights_array[4415:4384];      weights[647]=weights_array[4383:4352];      weights[648]=weights_array[4351:4320];      weights[649]=weights_array[4319:4288];      weights[650]=weights_array[4287:4256];      weights[651]=weights_array[4255:4224];      weights[652]=weights_array[4223:4192];      weights[653]=weights_array[4191:4160];      weights[654]=weights_array[4159:4128];      weights[655]=weights_array[4127:4096];      weights[656]=weights_array[4095:4064];      weights[657]=weights_array[4063:4032];      weights[658]=weights_array[4031:4000];      weights[659]=weights_array[3999:3968];      weights[660]=weights_array[3967:3936];      weights[661]=weights_array[3935:3904];      weights[662]=weights_array[3903:3872];      weights[663]=weights_array[3871:3840];      weights[664]=weights_array[3839:3808];      weights[665]=weights_array[3807:3776];      weights[666]=weights_array[3775:3744];      weights[667]=weights_array[3743:3712];      weights[668]=weights_array[3711:3680];      weights[669]=weights_array[3679:3648];      weights[670]=weights_array[3647:3616];      weights[671]=weights_array[3615:3584];      weights[672]=weights_array[3583:3552];      weights[673]=weights_array[3551:3520];      weights[674]=weights_array[3519:3488];      weights[675]=weights_array[3487:3456];      weights[676]=weights_array[3455:3424];      weights[677]=weights_array[3423:3392];      weights[678]=weights_array[3391:3360];      weights[679]=weights_array[3359:3328];      weights[680]=weights_array[3327:3296];      weights[681]=weights_array[3295:3264];      weights[682]=weights_array[3263:3232];      weights[683]=weights_array[3231:3200];      weights[684]=weights_array[3199:3168];      weights[685]=weights_array[3167:3136];      weights[686]=weights_array[3135:3104];      weights[687]=weights_array[3103:3072];      weights[688]=weights_array[3071:3040];      weights[689]=weights_array[3039:3008];      weights[690]=weights_array[3007:2976];      weights[691]=weights_array[2975:2944];      weights[692]=weights_array[2943:2912];      weights[693]=weights_array[2911:2880];      weights[694]=weights_array[2879:2848];      weights[695]=weights_array[2847:2816];      weights[696]=weights_array[2815:2784];      weights[697]=weights_array[2783:2752];      weights[698]=weights_array[2751:2720];      weights[699]=weights_array[2719:2688];      weights[700]=weights_array[2687:2656];      weights[701]=weights_array[2655:2624];      weights[702]=weights_array[2623:2592];      weights[703]=weights_array[2591:2560];      weights[704]=weights_array[2559:2528];      weights[705]=weights_array[2527:2496];      weights[706]=weights_array[2495:2464];      weights[707]=weights_array[2463:2432];      weights[708]=weights_array[2431:2400];      weights[709]=weights_array[2399:2368];      weights[710]=weights_array[2367:2336];      weights[711]=weights_array[2335:2304];      weights[712]=weights_array[2303:2272];      weights[713]=weights_array[2271:2240];      weights[714]=weights_array[2239:2208];      weights[715]=weights_array[2207:2176];      weights[716]=weights_array[2175:2144];      weights[717]=weights_array[2143:2112];      weights[718]=weights_array[2111:2080];      weights[719]=weights_array[2079:2048];      weights[720]=weights_array[2047:2016];      weights[721]=weights_array[2015:1984];      weights[722]=weights_array[1983:1952];      weights[723]=weights_array[1951:1920];      weights[724]=weights_array[1919:1888];      weights[725]=weights_array[1887:1856];      weights[726]=weights_array[1855:1824];      weights[727]=weights_array[1823:1792];      weights[728]=weights_array[1791:1760];      weights[729]=weights_array[1759:1728];      weights[730]=weights_array[1727:1696];      weights[731]=weights_array[1695:1664];      weights[732]=weights_array[1663:1632];      weights[733]=weights_array[1631:1600];      weights[734]=weights_array[1599:1568];      weights[735]=weights_array[1567:1536];      weights[736]=weights_array[1535:1504];      weights[737]=weights_array[1503:1472];      weights[738]=weights_array[1471:1440];      weights[739]=weights_array[1439:1408];      weights[740]=weights_array[1407:1376];      weights[741]=weights_array[1375:1344];      weights[742]=weights_array[1343:1312];      weights[743]=weights_array[1311:1280];      weights[744]=weights_array[1279:1248];      weights[745]=weights_array[1247:1216];      weights[746]=weights_array[1215:1184];      weights[747]=weights_array[1183:1152];      weights[748]=weights_array[1151:1120];      weights[749]=weights_array[1119:1088];      weights[750]=weights_array[1087:1056];      weights[751]=weights_array[1055:1024];      weights[752]=weights_array[1023:992];      weights[753]=weights_array[991:960];      weights[754]=weights_array[959:928];      weights[755]=weights_array[927:896];      weights[756]=weights_array[895:864];      weights[757]=weights_array[863:832];      weights[758]=weights_array[831:800];      weights[759]=weights_array[799:768];      weights[760]=weights_array[767:736];      weights[761]=weights_array[735:704];      weights[762]=weights_array[703:672];      weights[763]=weights_array[671:640];      weights[764]=weights_array[639:608];      weights[765]=weights_array[607:576];      weights[766]=weights_array[575:544];      weights[767]=weights_array[543:512];      weights[768]=weights_array[511:480];      weights[769]=weights_array[479:448];      weights[770]=weights_array[447:416];      weights[771]=weights_array[415:384];      weights[772]=weights_array[383:352];      weights[773]=weights_array[351:320];      weights[774]=weights_array[319:288];      weights[775]=weights_array[287:256];      weights[776]=weights_array[255:224];      weights[777]=weights_array[223:192];      weights[778]=weights_array[191:160];      weights[779]=weights_array[159:128];      weights[780]=weights_array[127:96];      weights[781]=weights_array[95:64];      weights[782]=weights_array[63:32];      weights[783]=weights_array[31:0];      
        // weights[4] = weights_array[31:0];
        // weights[3] = weights_array[63:32];
        // weights[2] = weights_array[95:64];
        // weights[1] = weights_array[127:96];
        // weights[0] = weights_array[159:128];

        //extract the initialization source address
source_addresses[0]=source_addresses_array[9407:9396];      source_addresses[1]=source_addresses_array[9395:9384];      source_addresses[2]=source_addresses_array[9383:9372];      source_addresses[3]=source_addresses_array[9371:9360];      source_addresses[4]=source_addresses_array[9359:9348];      source_addresses[5]=source_addresses_array[9347:9336];      source_addresses[6]=source_addresses_array[9335:9324];      source_addresses[7]=source_addresses_array[9323:9312];      source_addresses[8]=source_addresses_array[9311:9300];      source_addresses[9]=source_addresses_array[9299:9288];      source_addresses[10]=source_addresses_array[9287:9276];      source_addresses[11]=source_addresses_array[9275:9264];      source_addresses[12]=source_addresses_array[9263:9252];      source_addresses[13]=source_addresses_array[9251:9240];      source_addresses[14]=source_addresses_array[9239:9228];      source_addresses[15]=source_addresses_array[9227:9216];      source_addresses[16]=source_addresses_array[9215:9204];      source_addresses[17]=source_addresses_array[9203:9192];      source_addresses[18]=source_addresses_array[9191:9180];      source_addresses[19]=source_addresses_array[9179:9168];      source_addresses[20]=source_addresses_array[9167:9156];      source_addresses[21]=source_addresses_array[9155:9144];      source_addresses[22]=source_addresses_array[9143:9132];      source_addresses[23]=source_addresses_array[9131:9120];      source_addresses[24]=source_addresses_array[9119:9108];      source_addresses[25]=source_addresses_array[9107:9096];      source_addresses[26]=source_addresses_array[9095:9084];      source_addresses[27]=source_addresses_array[9083:9072];      source_addresses[28]=source_addresses_array[9071:9060];      source_addresses[29]=source_addresses_array[9059:9048];      source_addresses[30]=source_addresses_array[9047:9036];      source_addresses[31]=source_addresses_array[9035:9024];      source_addresses[32]=source_addresses_array[9023:9012];      source_addresses[33]=source_addresses_array[9011:9000];      source_addresses[34]=source_addresses_array[8999:8988];      source_addresses[35]=source_addresses_array[8987:8976];      source_addresses[36]=source_addresses_array[8975:8964];      source_addresses[37]=source_addresses_array[8963:8952];      source_addresses[38]=source_addresses_array[8951:8940];      source_addresses[39]=source_addresses_array[8939:8928];      source_addresses[40]=source_addresses_array[8927:8916];      source_addresses[41]=source_addresses_array[8915:8904];      source_addresses[42]=source_addresses_array[8903:8892];      source_addresses[43]=source_addresses_array[8891:8880];      source_addresses[44]=source_addresses_array[8879:8868];      source_addresses[45]=source_addresses_array[8867:8856];      source_addresses[46]=source_addresses_array[8855:8844];      source_addresses[47]=source_addresses_array[8843:8832];      source_addresses[48]=source_addresses_array[8831:8820];      source_addresses[49]=source_addresses_array[8819:8808];      source_addresses[50]=source_addresses_array[8807:8796];      source_addresses[51]=source_addresses_array[8795:8784];      source_addresses[52]=source_addresses_array[8783:8772];      source_addresses[53]=source_addresses_array[8771:8760];      source_addresses[54]=source_addresses_array[8759:8748];      source_addresses[55]=source_addresses_array[8747:8736];      source_addresses[56]=source_addresses_array[8735:8724];      source_addresses[57]=source_addresses_array[8723:8712];      source_addresses[58]=source_addresses_array[8711:8700];      source_addresses[59]=source_addresses_array[8699:8688];      source_addresses[60]=source_addresses_array[8687:8676];      source_addresses[61]=source_addresses_array[8675:8664];      source_addresses[62]=source_addresses_array[8663:8652];      source_addresses[63]=source_addresses_array[8651:8640];      source_addresses[64]=source_addresses_array[8639:8628];      source_addresses[65]=source_addresses_array[8627:8616];      source_addresses[66]=source_addresses_array[8615:8604];      source_addresses[67]=source_addresses_array[8603:8592];      source_addresses[68]=source_addresses_array[8591:8580];      source_addresses[69]=source_addresses_array[8579:8568];      source_addresses[70]=source_addresses_array[8567:8556];      source_addresses[71]=source_addresses_array[8555:8544];      source_addresses[72]=source_addresses_array[8543:8532];      source_addresses[73]=source_addresses_array[8531:8520];      source_addresses[74]=source_addresses_array[8519:8508];      source_addresses[75]=source_addresses_array[8507:8496];      source_addresses[76]=source_addresses_array[8495:8484];      source_addresses[77]=source_addresses_array[8483:8472];      source_addresses[78]=source_addresses_array[8471:8460];      source_addresses[79]=source_addresses_array[8459:8448];      source_addresses[80]=source_addresses_array[8447:8436];      source_addresses[81]=source_addresses_array[8435:8424];      source_addresses[82]=source_addresses_array[8423:8412];      source_addresses[83]=source_addresses_array[8411:8400];      source_addresses[84]=source_addresses_array[8399:8388];      source_addresses[85]=source_addresses_array[8387:8376];      source_addresses[86]=source_addresses_array[8375:8364];      source_addresses[87]=source_addresses_array[8363:8352];      source_addresses[88]=source_addresses_array[8351:8340];      source_addresses[89]=source_addresses_array[8339:8328];      source_addresses[90]=source_addresses_array[8327:8316];      source_addresses[91]=source_addresses_array[8315:8304];      source_addresses[92]=source_addresses_array[8303:8292];      source_addresses[93]=source_addresses_array[8291:8280];      source_addresses[94]=source_addresses_array[8279:8268];      source_addresses[95]=source_addresses_array[8267:8256];      source_addresses[96]=source_addresses_array[8255:8244];      source_addresses[97]=source_addresses_array[8243:8232];      source_addresses[98]=source_addresses_array[8231:8220];      source_addresses[99]=source_addresses_array[8219:8208];      source_addresses[100]=source_addresses_array[8207:8196];      source_addresses[101]=source_addresses_array[8195:8184];      source_addresses[102]=source_addresses_array[8183:8172];      source_addresses[103]=source_addresses_array[8171:8160];      source_addresses[104]=source_addresses_array[8159:8148];      source_addresses[105]=source_addresses_array[8147:8136];      source_addresses[106]=source_addresses_array[8135:8124];      source_addresses[107]=source_addresses_array[8123:8112];      source_addresses[108]=source_addresses_array[8111:8100];      source_addresses[109]=source_addresses_array[8099:8088];      source_addresses[110]=source_addresses_array[8087:8076];      source_addresses[111]=source_addresses_array[8075:8064];      source_addresses[112]=source_addresses_array[8063:8052];      source_addresses[113]=source_addresses_array[8051:8040];      source_addresses[114]=source_addresses_array[8039:8028];      source_addresses[115]=source_addresses_array[8027:8016];      source_addresses[116]=source_addresses_array[8015:8004];      source_addresses[117]=source_addresses_array[8003:7992];      source_addresses[118]=source_addresses_array[7991:7980];      source_addresses[119]=source_addresses_array[7979:7968];      source_addresses[120]=source_addresses_array[7967:7956];      source_addresses[121]=source_addresses_array[7955:7944];      source_addresses[122]=source_addresses_array[7943:7932];      source_addresses[123]=source_addresses_array[7931:7920];      source_addresses[124]=source_addresses_array[7919:7908];      source_addresses[125]=source_addresses_array[7907:7896];      source_addresses[126]=source_addresses_array[7895:7884];      source_addresses[127]=source_addresses_array[7883:7872];      source_addresses[128]=source_addresses_array[7871:7860];      source_addresses[129]=source_addresses_array[7859:7848];      source_addresses[130]=source_addresses_array[7847:7836];      source_addresses[131]=source_addresses_array[7835:7824];      source_addresses[132]=source_addresses_array[7823:7812];      source_addresses[133]=source_addresses_array[7811:7800];      source_addresses[134]=source_addresses_array[7799:7788];      source_addresses[135]=source_addresses_array[7787:7776];      source_addresses[136]=source_addresses_array[7775:7764];      source_addresses[137]=source_addresses_array[7763:7752];      source_addresses[138]=source_addresses_array[7751:7740];      source_addresses[139]=source_addresses_array[7739:7728];      source_addresses[140]=source_addresses_array[7727:7716];      source_addresses[141]=source_addresses_array[7715:7704];      source_addresses[142]=source_addresses_array[7703:7692];      source_addresses[143]=source_addresses_array[7691:7680];      source_addresses[144]=source_addresses_array[7679:7668];      source_addresses[145]=source_addresses_array[7667:7656];      source_addresses[146]=source_addresses_array[7655:7644];      source_addresses[147]=source_addresses_array[7643:7632];      source_addresses[148]=source_addresses_array[7631:7620];      source_addresses[149]=source_addresses_array[7619:7608];      source_addresses[150]=source_addresses_array[7607:7596];      source_addresses[151]=source_addresses_array[7595:7584];      source_addresses[152]=source_addresses_array[7583:7572];      source_addresses[153]=source_addresses_array[7571:7560];      source_addresses[154]=source_addresses_array[7559:7548];      source_addresses[155]=source_addresses_array[7547:7536];      source_addresses[156]=source_addresses_array[7535:7524];      source_addresses[157]=source_addresses_array[7523:7512];      source_addresses[158]=source_addresses_array[7511:7500];      source_addresses[159]=source_addresses_array[7499:7488];      source_addresses[160]=source_addresses_array[7487:7476];      source_addresses[161]=source_addresses_array[7475:7464];      source_addresses[162]=source_addresses_array[7463:7452];      source_addresses[163]=source_addresses_array[7451:7440];      source_addresses[164]=source_addresses_array[7439:7428];      source_addresses[165]=source_addresses_array[7427:7416];      source_addresses[166]=source_addresses_array[7415:7404];      source_addresses[167]=source_addresses_array[7403:7392];      source_addresses[168]=source_addresses_array[7391:7380];      source_addresses[169]=source_addresses_array[7379:7368];      source_addresses[170]=source_addresses_array[7367:7356];      source_addresses[171]=source_addresses_array[7355:7344];      source_addresses[172]=source_addresses_array[7343:7332];      source_addresses[173]=source_addresses_array[7331:7320];      source_addresses[174]=source_addresses_array[7319:7308];      source_addresses[175]=source_addresses_array[7307:7296];      source_addresses[176]=source_addresses_array[7295:7284];      source_addresses[177]=source_addresses_array[7283:7272];      source_addresses[178]=source_addresses_array[7271:7260];      source_addresses[179]=source_addresses_array[7259:7248];      source_addresses[180]=source_addresses_array[7247:7236];      source_addresses[181]=source_addresses_array[7235:7224];      source_addresses[182]=source_addresses_array[7223:7212];      source_addresses[183]=source_addresses_array[7211:7200];      source_addresses[184]=source_addresses_array[7199:7188];      source_addresses[185]=source_addresses_array[7187:7176];      source_addresses[186]=source_addresses_array[7175:7164];      source_addresses[187]=source_addresses_array[7163:7152];      source_addresses[188]=source_addresses_array[7151:7140];      source_addresses[189]=source_addresses_array[7139:7128];      source_addresses[190]=source_addresses_array[7127:7116];      source_addresses[191]=source_addresses_array[7115:7104];      source_addresses[192]=source_addresses_array[7103:7092];      source_addresses[193]=source_addresses_array[7091:7080];      source_addresses[194]=source_addresses_array[7079:7068];      source_addresses[195]=source_addresses_array[7067:7056];      source_addresses[196]=source_addresses_array[7055:7044];      source_addresses[197]=source_addresses_array[7043:7032];      source_addresses[198]=source_addresses_array[7031:7020];      source_addresses[199]=source_addresses_array[7019:7008];      source_addresses[200]=source_addresses_array[7007:6996];      source_addresses[201]=source_addresses_array[6995:6984];      source_addresses[202]=source_addresses_array[6983:6972];      source_addresses[203]=source_addresses_array[6971:6960];      source_addresses[204]=source_addresses_array[6959:6948];      source_addresses[205]=source_addresses_array[6947:6936];      source_addresses[206]=source_addresses_array[6935:6924];      source_addresses[207]=source_addresses_array[6923:6912];      source_addresses[208]=source_addresses_array[6911:6900];      source_addresses[209]=source_addresses_array[6899:6888];      source_addresses[210]=source_addresses_array[6887:6876];      source_addresses[211]=source_addresses_array[6875:6864];      source_addresses[212]=source_addresses_array[6863:6852];      source_addresses[213]=source_addresses_array[6851:6840];      source_addresses[214]=source_addresses_array[6839:6828];      source_addresses[215]=source_addresses_array[6827:6816];      source_addresses[216]=source_addresses_array[6815:6804];      source_addresses[217]=source_addresses_array[6803:6792];      source_addresses[218]=source_addresses_array[6791:6780];      source_addresses[219]=source_addresses_array[6779:6768];      source_addresses[220]=source_addresses_array[6767:6756];      source_addresses[221]=source_addresses_array[6755:6744];      source_addresses[222]=source_addresses_array[6743:6732];      source_addresses[223]=source_addresses_array[6731:6720];      source_addresses[224]=source_addresses_array[6719:6708];      source_addresses[225]=source_addresses_array[6707:6696];      source_addresses[226]=source_addresses_array[6695:6684];      source_addresses[227]=source_addresses_array[6683:6672];      source_addresses[228]=source_addresses_array[6671:6660];      source_addresses[229]=source_addresses_array[6659:6648];      source_addresses[230]=source_addresses_array[6647:6636];      source_addresses[231]=source_addresses_array[6635:6624];      source_addresses[232]=source_addresses_array[6623:6612];      source_addresses[233]=source_addresses_array[6611:6600];      source_addresses[234]=source_addresses_array[6599:6588];      source_addresses[235]=source_addresses_array[6587:6576];      source_addresses[236]=source_addresses_array[6575:6564];      source_addresses[237]=source_addresses_array[6563:6552];      source_addresses[238]=source_addresses_array[6551:6540];      source_addresses[239]=source_addresses_array[6539:6528];      source_addresses[240]=source_addresses_array[6527:6516];      source_addresses[241]=source_addresses_array[6515:6504];      source_addresses[242]=source_addresses_array[6503:6492];      source_addresses[243]=source_addresses_array[6491:6480];      source_addresses[244]=source_addresses_array[6479:6468];      source_addresses[245]=source_addresses_array[6467:6456];      source_addresses[246]=source_addresses_array[6455:6444];      source_addresses[247]=source_addresses_array[6443:6432];      source_addresses[248]=source_addresses_array[6431:6420];      source_addresses[249]=source_addresses_array[6419:6408];      source_addresses[250]=source_addresses_array[6407:6396];      source_addresses[251]=source_addresses_array[6395:6384];      source_addresses[252]=source_addresses_array[6383:6372];      source_addresses[253]=source_addresses_array[6371:6360];      source_addresses[254]=source_addresses_array[6359:6348];      source_addresses[255]=source_addresses_array[6347:6336];      source_addresses[256]=source_addresses_array[6335:6324];      source_addresses[257]=source_addresses_array[6323:6312];      source_addresses[258]=source_addresses_array[6311:6300];      source_addresses[259]=source_addresses_array[6299:6288];      source_addresses[260]=source_addresses_array[6287:6276];      source_addresses[261]=source_addresses_array[6275:6264];      source_addresses[262]=source_addresses_array[6263:6252];      source_addresses[263]=source_addresses_array[6251:6240];      source_addresses[264]=source_addresses_array[6239:6228];      source_addresses[265]=source_addresses_array[6227:6216];      source_addresses[266]=source_addresses_array[6215:6204];      source_addresses[267]=source_addresses_array[6203:6192];      source_addresses[268]=source_addresses_array[6191:6180];      source_addresses[269]=source_addresses_array[6179:6168];      source_addresses[270]=source_addresses_array[6167:6156];      source_addresses[271]=source_addresses_array[6155:6144];      source_addresses[272]=source_addresses_array[6143:6132];      source_addresses[273]=source_addresses_array[6131:6120];      source_addresses[274]=source_addresses_array[6119:6108];      source_addresses[275]=source_addresses_array[6107:6096];      source_addresses[276]=source_addresses_array[6095:6084];      source_addresses[277]=source_addresses_array[6083:6072];      source_addresses[278]=source_addresses_array[6071:6060];      source_addresses[279]=source_addresses_array[6059:6048];      source_addresses[280]=source_addresses_array[6047:6036];      source_addresses[281]=source_addresses_array[6035:6024];      source_addresses[282]=source_addresses_array[6023:6012];      source_addresses[283]=source_addresses_array[6011:6000];      source_addresses[284]=source_addresses_array[5999:5988];      source_addresses[285]=source_addresses_array[5987:5976];      source_addresses[286]=source_addresses_array[5975:5964];      source_addresses[287]=source_addresses_array[5963:5952];      source_addresses[288]=source_addresses_array[5951:5940];      source_addresses[289]=source_addresses_array[5939:5928];      source_addresses[290]=source_addresses_array[5927:5916];      source_addresses[291]=source_addresses_array[5915:5904];      source_addresses[292]=source_addresses_array[5903:5892];      source_addresses[293]=source_addresses_array[5891:5880];      source_addresses[294]=source_addresses_array[5879:5868];      source_addresses[295]=source_addresses_array[5867:5856];      source_addresses[296]=source_addresses_array[5855:5844];      source_addresses[297]=source_addresses_array[5843:5832];      source_addresses[298]=source_addresses_array[5831:5820];      source_addresses[299]=source_addresses_array[5819:5808];      source_addresses[300]=source_addresses_array[5807:5796];      source_addresses[301]=source_addresses_array[5795:5784];      source_addresses[302]=source_addresses_array[5783:5772];      source_addresses[303]=source_addresses_array[5771:5760];      source_addresses[304]=source_addresses_array[5759:5748];      source_addresses[305]=source_addresses_array[5747:5736];      source_addresses[306]=source_addresses_array[5735:5724];      source_addresses[307]=source_addresses_array[5723:5712];      source_addresses[308]=source_addresses_array[5711:5700];      source_addresses[309]=source_addresses_array[5699:5688];      source_addresses[310]=source_addresses_array[5687:5676];      source_addresses[311]=source_addresses_array[5675:5664];      source_addresses[312]=source_addresses_array[5663:5652];      source_addresses[313]=source_addresses_array[5651:5640];      source_addresses[314]=source_addresses_array[5639:5628];      source_addresses[315]=source_addresses_array[5627:5616];      source_addresses[316]=source_addresses_array[5615:5604];      source_addresses[317]=source_addresses_array[5603:5592];      source_addresses[318]=source_addresses_array[5591:5580];      source_addresses[319]=source_addresses_array[5579:5568];      source_addresses[320]=source_addresses_array[5567:5556];      source_addresses[321]=source_addresses_array[5555:5544];      source_addresses[322]=source_addresses_array[5543:5532];      source_addresses[323]=source_addresses_array[5531:5520];      source_addresses[324]=source_addresses_array[5519:5508];      source_addresses[325]=source_addresses_array[5507:5496];      source_addresses[326]=source_addresses_array[5495:5484];      source_addresses[327]=source_addresses_array[5483:5472];      source_addresses[328]=source_addresses_array[5471:5460];      source_addresses[329]=source_addresses_array[5459:5448];      source_addresses[330]=source_addresses_array[5447:5436];      source_addresses[331]=source_addresses_array[5435:5424];      source_addresses[332]=source_addresses_array[5423:5412];      source_addresses[333]=source_addresses_array[5411:5400];      source_addresses[334]=source_addresses_array[5399:5388];      source_addresses[335]=source_addresses_array[5387:5376];      source_addresses[336]=source_addresses_array[5375:5364];      source_addresses[337]=source_addresses_array[5363:5352];      source_addresses[338]=source_addresses_array[5351:5340];      source_addresses[339]=source_addresses_array[5339:5328];      source_addresses[340]=source_addresses_array[5327:5316];      source_addresses[341]=source_addresses_array[5315:5304];      source_addresses[342]=source_addresses_array[5303:5292];      source_addresses[343]=source_addresses_array[5291:5280];      source_addresses[344]=source_addresses_array[5279:5268];      source_addresses[345]=source_addresses_array[5267:5256];      source_addresses[346]=source_addresses_array[5255:5244];      source_addresses[347]=source_addresses_array[5243:5232];      source_addresses[348]=source_addresses_array[5231:5220];      source_addresses[349]=source_addresses_array[5219:5208];      source_addresses[350]=source_addresses_array[5207:5196];      source_addresses[351]=source_addresses_array[5195:5184];      source_addresses[352]=source_addresses_array[5183:5172];      source_addresses[353]=source_addresses_array[5171:5160];      source_addresses[354]=source_addresses_array[5159:5148];      source_addresses[355]=source_addresses_array[5147:5136];      source_addresses[356]=source_addresses_array[5135:5124];      source_addresses[357]=source_addresses_array[5123:5112];      source_addresses[358]=source_addresses_array[5111:5100];      source_addresses[359]=source_addresses_array[5099:5088];      source_addresses[360]=source_addresses_array[5087:5076];      source_addresses[361]=source_addresses_array[5075:5064];      source_addresses[362]=source_addresses_array[5063:5052];      source_addresses[363]=source_addresses_array[5051:5040];      source_addresses[364]=source_addresses_array[5039:5028];      source_addresses[365]=source_addresses_array[5027:5016];      source_addresses[366]=source_addresses_array[5015:5004];      source_addresses[367]=source_addresses_array[5003:4992];      source_addresses[368]=source_addresses_array[4991:4980];      source_addresses[369]=source_addresses_array[4979:4968];      source_addresses[370]=source_addresses_array[4967:4956];      source_addresses[371]=source_addresses_array[4955:4944];      source_addresses[372]=source_addresses_array[4943:4932];      source_addresses[373]=source_addresses_array[4931:4920];      source_addresses[374]=source_addresses_array[4919:4908];      source_addresses[375]=source_addresses_array[4907:4896];      source_addresses[376]=source_addresses_array[4895:4884];      source_addresses[377]=source_addresses_array[4883:4872];      source_addresses[378]=source_addresses_array[4871:4860];      source_addresses[379]=source_addresses_array[4859:4848];      source_addresses[380]=source_addresses_array[4847:4836];      source_addresses[381]=source_addresses_array[4835:4824];      source_addresses[382]=source_addresses_array[4823:4812];      source_addresses[383]=source_addresses_array[4811:4800];      source_addresses[384]=source_addresses_array[4799:4788];      source_addresses[385]=source_addresses_array[4787:4776];      source_addresses[386]=source_addresses_array[4775:4764];      source_addresses[387]=source_addresses_array[4763:4752];      source_addresses[388]=source_addresses_array[4751:4740];      source_addresses[389]=source_addresses_array[4739:4728];      source_addresses[390]=source_addresses_array[4727:4716];      source_addresses[391]=source_addresses_array[4715:4704];      source_addresses[392]=source_addresses_array[4703:4692];      source_addresses[393]=source_addresses_array[4691:4680];      source_addresses[394]=source_addresses_array[4679:4668];      source_addresses[395]=source_addresses_array[4667:4656];      source_addresses[396]=source_addresses_array[4655:4644];      source_addresses[397]=source_addresses_array[4643:4632];      source_addresses[398]=source_addresses_array[4631:4620];      source_addresses[399]=source_addresses_array[4619:4608];      source_addresses[400]=source_addresses_array[4607:4596];      source_addresses[401]=source_addresses_array[4595:4584];      source_addresses[402]=source_addresses_array[4583:4572];      source_addresses[403]=source_addresses_array[4571:4560];      source_addresses[404]=source_addresses_array[4559:4548];      source_addresses[405]=source_addresses_array[4547:4536];      source_addresses[406]=source_addresses_array[4535:4524];      source_addresses[407]=source_addresses_array[4523:4512];      source_addresses[408]=source_addresses_array[4511:4500];      source_addresses[409]=source_addresses_array[4499:4488];      source_addresses[410]=source_addresses_array[4487:4476];      source_addresses[411]=source_addresses_array[4475:4464];      source_addresses[412]=source_addresses_array[4463:4452];      source_addresses[413]=source_addresses_array[4451:4440];      source_addresses[414]=source_addresses_array[4439:4428];      source_addresses[415]=source_addresses_array[4427:4416];      source_addresses[416]=source_addresses_array[4415:4404];      source_addresses[417]=source_addresses_array[4403:4392];      source_addresses[418]=source_addresses_array[4391:4380];      source_addresses[419]=source_addresses_array[4379:4368];      source_addresses[420]=source_addresses_array[4367:4356];      source_addresses[421]=source_addresses_array[4355:4344];      source_addresses[422]=source_addresses_array[4343:4332];      source_addresses[423]=source_addresses_array[4331:4320];      source_addresses[424]=source_addresses_array[4319:4308];      source_addresses[425]=source_addresses_array[4307:4296];      source_addresses[426]=source_addresses_array[4295:4284];      source_addresses[427]=source_addresses_array[4283:4272];      source_addresses[428]=source_addresses_array[4271:4260];      source_addresses[429]=source_addresses_array[4259:4248];      source_addresses[430]=source_addresses_array[4247:4236];      source_addresses[431]=source_addresses_array[4235:4224];      source_addresses[432]=source_addresses_array[4223:4212];      source_addresses[433]=source_addresses_array[4211:4200];      source_addresses[434]=source_addresses_array[4199:4188];      source_addresses[435]=source_addresses_array[4187:4176];      source_addresses[436]=source_addresses_array[4175:4164];      source_addresses[437]=source_addresses_array[4163:4152];      source_addresses[438]=source_addresses_array[4151:4140];      source_addresses[439]=source_addresses_array[4139:4128];      source_addresses[440]=source_addresses_array[4127:4116];      source_addresses[441]=source_addresses_array[4115:4104];      source_addresses[442]=source_addresses_array[4103:4092];      source_addresses[443]=source_addresses_array[4091:4080];      source_addresses[444]=source_addresses_array[4079:4068];      source_addresses[445]=source_addresses_array[4067:4056];      source_addresses[446]=source_addresses_array[4055:4044];      source_addresses[447]=source_addresses_array[4043:4032];      source_addresses[448]=source_addresses_array[4031:4020];      source_addresses[449]=source_addresses_array[4019:4008];      source_addresses[450]=source_addresses_array[4007:3996];      source_addresses[451]=source_addresses_array[3995:3984];      source_addresses[452]=source_addresses_array[3983:3972];      source_addresses[453]=source_addresses_array[3971:3960];      source_addresses[454]=source_addresses_array[3959:3948];      source_addresses[455]=source_addresses_array[3947:3936];      source_addresses[456]=source_addresses_array[3935:3924];      source_addresses[457]=source_addresses_array[3923:3912];      source_addresses[458]=source_addresses_array[3911:3900];      source_addresses[459]=source_addresses_array[3899:3888];      source_addresses[460]=source_addresses_array[3887:3876];      source_addresses[461]=source_addresses_array[3875:3864];      source_addresses[462]=source_addresses_array[3863:3852];      source_addresses[463]=source_addresses_array[3851:3840];      source_addresses[464]=source_addresses_array[3839:3828];      source_addresses[465]=source_addresses_array[3827:3816];      source_addresses[466]=source_addresses_array[3815:3804];      source_addresses[467]=source_addresses_array[3803:3792];      source_addresses[468]=source_addresses_array[3791:3780];      source_addresses[469]=source_addresses_array[3779:3768];      source_addresses[470]=source_addresses_array[3767:3756];      source_addresses[471]=source_addresses_array[3755:3744];      source_addresses[472]=source_addresses_array[3743:3732];      source_addresses[473]=source_addresses_array[3731:3720];      source_addresses[474]=source_addresses_array[3719:3708];      source_addresses[475]=source_addresses_array[3707:3696];      source_addresses[476]=source_addresses_array[3695:3684];      source_addresses[477]=source_addresses_array[3683:3672];      source_addresses[478]=source_addresses_array[3671:3660];      source_addresses[479]=source_addresses_array[3659:3648];      source_addresses[480]=source_addresses_array[3647:3636];      source_addresses[481]=source_addresses_array[3635:3624];      source_addresses[482]=source_addresses_array[3623:3612];      source_addresses[483]=source_addresses_array[3611:3600];      source_addresses[484]=source_addresses_array[3599:3588];      source_addresses[485]=source_addresses_array[3587:3576];      source_addresses[486]=source_addresses_array[3575:3564];      source_addresses[487]=source_addresses_array[3563:3552];      source_addresses[488]=source_addresses_array[3551:3540];      source_addresses[489]=source_addresses_array[3539:3528];      source_addresses[490]=source_addresses_array[3527:3516];      source_addresses[491]=source_addresses_array[3515:3504];      source_addresses[492]=source_addresses_array[3503:3492];      source_addresses[493]=source_addresses_array[3491:3480];      source_addresses[494]=source_addresses_array[3479:3468];      source_addresses[495]=source_addresses_array[3467:3456];      source_addresses[496]=source_addresses_array[3455:3444];      source_addresses[497]=source_addresses_array[3443:3432];      source_addresses[498]=source_addresses_array[3431:3420];      source_addresses[499]=source_addresses_array[3419:3408];      source_addresses[500]=source_addresses_array[3407:3396];      source_addresses[501]=source_addresses_array[3395:3384];      source_addresses[502]=source_addresses_array[3383:3372];      source_addresses[503]=source_addresses_array[3371:3360];      source_addresses[504]=source_addresses_array[3359:3348];      source_addresses[505]=source_addresses_array[3347:3336];      source_addresses[506]=source_addresses_array[3335:3324];      source_addresses[507]=source_addresses_array[3323:3312];      source_addresses[508]=source_addresses_array[3311:3300];      source_addresses[509]=source_addresses_array[3299:3288];      source_addresses[510]=source_addresses_array[3287:3276];      source_addresses[511]=source_addresses_array[3275:3264];      source_addresses[512]=source_addresses_array[3263:3252];      source_addresses[513]=source_addresses_array[3251:3240];      source_addresses[514]=source_addresses_array[3239:3228];      source_addresses[515]=source_addresses_array[3227:3216];      source_addresses[516]=source_addresses_array[3215:3204];      source_addresses[517]=source_addresses_array[3203:3192];      source_addresses[518]=source_addresses_array[3191:3180];      source_addresses[519]=source_addresses_array[3179:3168];      source_addresses[520]=source_addresses_array[3167:3156];      source_addresses[521]=source_addresses_array[3155:3144];      source_addresses[522]=source_addresses_array[3143:3132];      source_addresses[523]=source_addresses_array[3131:3120];      source_addresses[524]=source_addresses_array[3119:3108];      source_addresses[525]=source_addresses_array[3107:3096];      source_addresses[526]=source_addresses_array[3095:3084];      source_addresses[527]=source_addresses_array[3083:3072];      source_addresses[528]=source_addresses_array[3071:3060];      source_addresses[529]=source_addresses_array[3059:3048];      source_addresses[530]=source_addresses_array[3047:3036];      source_addresses[531]=source_addresses_array[3035:3024];      source_addresses[532]=source_addresses_array[3023:3012];      source_addresses[533]=source_addresses_array[3011:3000];      source_addresses[534]=source_addresses_array[2999:2988];      source_addresses[535]=source_addresses_array[2987:2976];      source_addresses[536]=source_addresses_array[2975:2964];      source_addresses[537]=source_addresses_array[2963:2952];      source_addresses[538]=source_addresses_array[2951:2940];      source_addresses[539]=source_addresses_array[2939:2928];      source_addresses[540]=source_addresses_array[2927:2916];      source_addresses[541]=source_addresses_array[2915:2904];      source_addresses[542]=source_addresses_array[2903:2892];      source_addresses[543]=source_addresses_array[2891:2880];      source_addresses[544]=source_addresses_array[2879:2868];      source_addresses[545]=source_addresses_array[2867:2856];      source_addresses[546]=source_addresses_array[2855:2844];      source_addresses[547]=source_addresses_array[2843:2832];      source_addresses[548]=source_addresses_array[2831:2820];      source_addresses[549]=source_addresses_array[2819:2808];      source_addresses[550]=source_addresses_array[2807:2796];      source_addresses[551]=source_addresses_array[2795:2784];      source_addresses[552]=source_addresses_array[2783:2772];      source_addresses[553]=source_addresses_array[2771:2760];      source_addresses[554]=source_addresses_array[2759:2748];      source_addresses[555]=source_addresses_array[2747:2736];      source_addresses[556]=source_addresses_array[2735:2724];      source_addresses[557]=source_addresses_array[2723:2712];      source_addresses[558]=source_addresses_array[2711:2700];      source_addresses[559]=source_addresses_array[2699:2688];      source_addresses[560]=source_addresses_array[2687:2676];      source_addresses[561]=source_addresses_array[2675:2664];      source_addresses[562]=source_addresses_array[2663:2652];      source_addresses[563]=source_addresses_array[2651:2640];      source_addresses[564]=source_addresses_array[2639:2628];      source_addresses[565]=source_addresses_array[2627:2616];      source_addresses[566]=source_addresses_array[2615:2604];      source_addresses[567]=source_addresses_array[2603:2592];      source_addresses[568]=source_addresses_array[2591:2580];      source_addresses[569]=source_addresses_array[2579:2568];      source_addresses[570]=source_addresses_array[2567:2556];      source_addresses[571]=source_addresses_array[2555:2544];      source_addresses[572]=source_addresses_array[2543:2532];      source_addresses[573]=source_addresses_array[2531:2520];      source_addresses[574]=source_addresses_array[2519:2508];      source_addresses[575]=source_addresses_array[2507:2496];      source_addresses[576]=source_addresses_array[2495:2484];      source_addresses[577]=source_addresses_array[2483:2472];      source_addresses[578]=source_addresses_array[2471:2460];      source_addresses[579]=source_addresses_array[2459:2448];      source_addresses[580]=source_addresses_array[2447:2436];      source_addresses[581]=source_addresses_array[2435:2424];      source_addresses[582]=source_addresses_array[2423:2412];      source_addresses[583]=source_addresses_array[2411:2400];      source_addresses[584]=source_addresses_array[2399:2388];      source_addresses[585]=source_addresses_array[2387:2376];      source_addresses[586]=source_addresses_array[2375:2364];      source_addresses[587]=source_addresses_array[2363:2352];      source_addresses[588]=source_addresses_array[2351:2340];      source_addresses[589]=source_addresses_array[2339:2328];      source_addresses[590]=source_addresses_array[2327:2316];      source_addresses[591]=source_addresses_array[2315:2304];      source_addresses[592]=source_addresses_array[2303:2292];      source_addresses[593]=source_addresses_array[2291:2280];      source_addresses[594]=source_addresses_array[2279:2268];      source_addresses[595]=source_addresses_array[2267:2256];      source_addresses[596]=source_addresses_array[2255:2244];      source_addresses[597]=source_addresses_array[2243:2232];      source_addresses[598]=source_addresses_array[2231:2220];      source_addresses[599]=source_addresses_array[2219:2208];      source_addresses[600]=source_addresses_array[2207:2196];      source_addresses[601]=source_addresses_array[2195:2184];      source_addresses[602]=source_addresses_array[2183:2172];      source_addresses[603]=source_addresses_array[2171:2160];      source_addresses[604]=source_addresses_array[2159:2148];      source_addresses[605]=source_addresses_array[2147:2136];      source_addresses[606]=source_addresses_array[2135:2124];      source_addresses[607]=source_addresses_array[2123:2112];      source_addresses[608]=source_addresses_array[2111:2100];      source_addresses[609]=source_addresses_array[2099:2088];      source_addresses[610]=source_addresses_array[2087:2076];      source_addresses[611]=source_addresses_array[2075:2064];      source_addresses[612]=source_addresses_array[2063:2052];      source_addresses[613]=source_addresses_array[2051:2040];      source_addresses[614]=source_addresses_array[2039:2028];      source_addresses[615]=source_addresses_array[2027:2016];      source_addresses[616]=source_addresses_array[2015:2004];      source_addresses[617]=source_addresses_array[2003:1992];      source_addresses[618]=source_addresses_array[1991:1980];      source_addresses[619]=source_addresses_array[1979:1968];      source_addresses[620]=source_addresses_array[1967:1956];      source_addresses[621]=source_addresses_array[1955:1944];      source_addresses[622]=source_addresses_array[1943:1932];      source_addresses[623]=source_addresses_array[1931:1920];      source_addresses[624]=source_addresses_array[1919:1908];      source_addresses[625]=source_addresses_array[1907:1896];      source_addresses[626]=source_addresses_array[1895:1884];      source_addresses[627]=source_addresses_array[1883:1872];      source_addresses[628]=source_addresses_array[1871:1860];      source_addresses[629]=source_addresses_array[1859:1848];      source_addresses[630]=source_addresses_array[1847:1836];      source_addresses[631]=source_addresses_array[1835:1824];      source_addresses[632]=source_addresses_array[1823:1812];      source_addresses[633]=source_addresses_array[1811:1800];      source_addresses[634]=source_addresses_array[1799:1788];      source_addresses[635]=source_addresses_array[1787:1776];      source_addresses[636]=source_addresses_array[1775:1764];      source_addresses[637]=source_addresses_array[1763:1752];      source_addresses[638]=source_addresses_array[1751:1740];      source_addresses[639]=source_addresses_array[1739:1728];      source_addresses[640]=source_addresses_array[1727:1716];      source_addresses[641]=source_addresses_array[1715:1704];      source_addresses[642]=source_addresses_array[1703:1692];      source_addresses[643]=source_addresses_array[1691:1680];      source_addresses[644]=source_addresses_array[1679:1668];      source_addresses[645]=source_addresses_array[1667:1656];      source_addresses[646]=source_addresses_array[1655:1644];      source_addresses[647]=source_addresses_array[1643:1632];      source_addresses[648]=source_addresses_array[1631:1620];      source_addresses[649]=source_addresses_array[1619:1608];      source_addresses[650]=source_addresses_array[1607:1596];      source_addresses[651]=source_addresses_array[1595:1584];      source_addresses[652]=source_addresses_array[1583:1572];      source_addresses[653]=source_addresses_array[1571:1560];      source_addresses[654]=source_addresses_array[1559:1548];      source_addresses[655]=source_addresses_array[1547:1536];      source_addresses[656]=source_addresses_array[1535:1524];      source_addresses[657]=source_addresses_array[1523:1512];      source_addresses[658]=source_addresses_array[1511:1500];      source_addresses[659]=source_addresses_array[1499:1488];      source_addresses[660]=source_addresses_array[1487:1476];      source_addresses[661]=source_addresses_array[1475:1464];      source_addresses[662]=source_addresses_array[1463:1452];      source_addresses[663]=source_addresses_array[1451:1440];      source_addresses[664]=source_addresses_array[1439:1428];      source_addresses[665]=source_addresses_array[1427:1416];      source_addresses[666]=source_addresses_array[1415:1404];      source_addresses[667]=source_addresses_array[1403:1392];      source_addresses[668]=source_addresses_array[1391:1380];      source_addresses[669]=source_addresses_array[1379:1368];      source_addresses[670]=source_addresses_array[1367:1356];      source_addresses[671]=source_addresses_array[1355:1344];      source_addresses[672]=source_addresses_array[1343:1332];      source_addresses[673]=source_addresses_array[1331:1320];      source_addresses[674]=source_addresses_array[1319:1308];      source_addresses[675]=source_addresses_array[1307:1296];      source_addresses[676]=source_addresses_array[1295:1284];      source_addresses[677]=source_addresses_array[1283:1272];      source_addresses[678]=source_addresses_array[1271:1260];      source_addresses[679]=source_addresses_array[1259:1248];      source_addresses[680]=source_addresses_array[1247:1236];      source_addresses[681]=source_addresses_array[1235:1224];      source_addresses[682]=source_addresses_array[1223:1212];      source_addresses[683]=source_addresses_array[1211:1200];      source_addresses[684]=source_addresses_array[1199:1188];      source_addresses[685]=source_addresses_array[1187:1176];      source_addresses[686]=source_addresses_array[1175:1164];      source_addresses[687]=source_addresses_array[1163:1152];      source_addresses[688]=source_addresses_array[1151:1140];      source_addresses[689]=source_addresses_array[1139:1128];      source_addresses[690]=source_addresses_array[1127:1116];      source_addresses[691]=source_addresses_array[1115:1104];      source_addresses[692]=source_addresses_array[1103:1092];      source_addresses[693]=source_addresses_array[1091:1080];      source_addresses[694]=source_addresses_array[1079:1068];      source_addresses[695]=source_addresses_array[1067:1056];      source_addresses[696]=source_addresses_array[1055:1044];      source_addresses[697]=source_addresses_array[1043:1032];      source_addresses[698]=source_addresses_array[1031:1020];      source_addresses[699]=source_addresses_array[1019:1008];      source_addresses[700]=source_addresses_array[1007:996];      source_addresses[701]=source_addresses_array[995:984];      source_addresses[702]=source_addresses_array[983:972];      source_addresses[703]=source_addresses_array[971:960];      source_addresses[704]=source_addresses_array[959:948];      source_addresses[705]=source_addresses_array[947:936];      source_addresses[706]=source_addresses_array[935:924];      source_addresses[707]=source_addresses_array[923:912];      source_addresses[708]=source_addresses_array[911:900];      source_addresses[709]=source_addresses_array[899:888];      source_addresses[710]=source_addresses_array[887:876];      source_addresses[711]=source_addresses_array[875:864];      source_addresses[712]=source_addresses_array[863:852];      source_addresses[713]=source_addresses_array[851:840];      source_addresses[714]=source_addresses_array[839:828];      source_addresses[715]=source_addresses_array[827:816];      source_addresses[716]=source_addresses_array[815:804];      source_addresses[717]=source_addresses_array[803:792];      source_addresses[718]=source_addresses_array[791:780];      source_addresses[719]=source_addresses_array[779:768];      source_addresses[720]=source_addresses_array[767:756];      source_addresses[721]=source_addresses_array[755:744];      source_addresses[722]=source_addresses_array[743:732];      source_addresses[723]=source_addresses_array[731:720];      source_addresses[724]=source_addresses_array[719:708];      source_addresses[725]=source_addresses_array[707:696];      source_addresses[726]=source_addresses_array[695:684];      source_addresses[727]=source_addresses_array[683:672];      source_addresses[728]=source_addresses_array[671:660];      source_addresses[729]=source_addresses_array[659:648];      source_addresses[730]=source_addresses_array[647:636];      source_addresses[731]=source_addresses_array[635:624];      source_addresses[732]=source_addresses_array[623:612];      source_addresses[733]=source_addresses_array[611:600];      source_addresses[734]=source_addresses_array[599:588];      source_addresses[735]=source_addresses_array[587:576];      source_addresses[736]=source_addresses_array[575:564];      source_addresses[737]=source_addresses_array[563:552];      source_addresses[738]=source_addresses_array[551:540];      source_addresses[739]=source_addresses_array[539:528];      source_addresses[740]=source_addresses_array[527:516];      source_addresses[741]=source_addresses_array[515:504];      source_addresses[742]=source_addresses_array[503:492];      source_addresses[743]=source_addresses_array[491:480];      source_addresses[744]=source_addresses_array[479:468];      source_addresses[745]=source_addresses_array[467:456];      source_addresses[746]=source_addresses_array[455:444];      source_addresses[747]=source_addresses_array[443:432];      source_addresses[748]=source_addresses_array[431:420];      source_addresses[749]=source_addresses_array[419:408];      source_addresses[750]=source_addresses_array[407:396];      source_addresses[751]=source_addresses_array[395:384];      source_addresses[752]=source_addresses_array[383:372];      source_addresses[753]=source_addresses_array[371:360];      source_addresses[754]=source_addresses_array[359:348];      source_addresses[755]=source_addresses_array[347:336];      source_addresses[756]=source_addresses_array[335:324];      source_addresses[757]=source_addresses_array[323:312];      source_addresses[758]=source_addresses_array[311:300];      source_addresses[759]=source_addresses_array[299:288];      source_addresses[760]=source_addresses_array[287:276];      source_addresses[761]=source_addresses_array[275:264];      source_addresses[762]=source_addresses_array[263:252];      source_addresses[763]=source_addresses_array[251:240];      source_addresses[764]=source_addresses_array[239:228];      source_addresses[765]=source_addresses_array[227:216];      source_addresses[766]=source_addresses_array[215:204];      source_addresses[767]=source_addresses_array[203:192];      source_addresses[768]=source_addresses_array[191:180];      source_addresses[769]=source_addresses_array[179:168];      source_addresses[770]=source_addresses_array[167:156];      source_addresses[771]=source_addresses_array[155:144];      source_addresses[772]=source_addresses_array[143:132];      source_addresses[773]=source_addresses_array[131:120];      source_addresses[774]=source_addresses_array[119:108];      source_addresses[775]=source_addresses_array[107:96];      source_addresses[776]=source_addresses_array[95:84];      source_addresses[777]=source_addresses_array[83:72];      source_addresses[778]=source_addresses_array[71:60];      source_addresses[779]=source_addresses_array[59:48];      source_addresses[780]=source_addresses_array[47:36];      source_addresses[781]=source_addresses_array[35:24];      source_addresses[782]=source_addresses_array[23:12];      source_addresses[783]=source_addresses_array[11:0];      
        // //break up the source adddresses
        // source_addresses[4] = source_addresses_array[11:0];
        // source_addresses[3] = source_addresses_array[23:12];
        // source_addresses[2] = source_addresses_array[35:24];
        // source_addresses[1] = source_addresses_array[47:36];
        // source_addresses[0] = source_addresses_array[59:48];
    end

    //when a spike/source address comes in get index and mark the incoming spike array
    always @(source_address) begin

        //get index by going through the source addresses
        break = 1'b0;
        for(i=0; i<number_of_connections; i=i+1) begin
            if (source_addresses[i] == source_address) begin
                index = i;
            end
        end

        incoming_spikes[index] = 1'b1;      //record the incoming spike
    end

    //when clear signal comes reset read the icnoming spike array and reset it
    always @(clear) begin
        case(clear)
            1'b1: begin
                for(i=0; i<number_of_connections; i=i+1) begin      //reset the incoming spikes array
                    spikes[i] = incoming_spikes[i];     //store the incoming spikes
                    incoming_spikes[i] = 1'b0;
                end

                accumulated_weight = 32'd0;     //set accumulated value to 0
                considered_weight = 32'd0;      //weight addition is zero

                //at the begining of the timestep accumulate weights and send to the potential adder unit
                for(i=0; i<number_of_connections; i=i+1) begin
                    if(spikes[i] == 1'b1) begin
                        #1
                        considered_weight <= weights[i];         
                        accumulated_weight <= added_weight;
                    end
                end
            end
        endcase
    end

    //added weight
    always @(added_weight) begin
        mult_output = added_weight;
    end


    initial begin
        //set incoming spikes array to zeros
        for(i=0; i<number_of_connections; i=i+1) begin      
            spikes[i] = 1'b0;    
            incoming_spikes[i] = 1'b0;
        end
    end


    // reg [127:0] mask;           //mask varibale to mask the weight that needs to be added
    // reg [127:0] mult_ans;       //weight answer after masking
    // reg [127:0] weight;         //4 weights at once
    // // For floating point addition
    // wire excpetion1, excpetion2, exception3;
    // wire [31:0] add_val1, add_val2, add_val3;

    //at the beginning of a timestep

    // always @(posedge CLK) begin 
    //     case (spike_in) 
    //         4'd0:   mult_output = 32'b0;                  // No spikes in any of the 4 branches.
    //         4'd1: begin
    //             mask = 128'b0;
    //             mask[31:0] = 32'd4294967295;   
    //             mult_ans = weight & mask; 
    //         end
    //         4'd2: begin
    //             mask = 128'b0;
    //             mask[63:32] = 32'd4294967295;   
    //             mult_ans = weight & mask; 
    //         end
    //         4'd3: begin
    //             mask = 128'b0;
    //             mask[63:0] = 32'd4294967295;   
    //             mult_ans = weight & mask; 
    //         end
    //         4'd4: begin
    //             mask = 128'b0;
    //             mask[95:64] = 32'd4294967295;   
    //             mult_ans = weight & mask; 
    //         end
    //         4'd5: begin
    //             mask = 128'b0;
    //             mask[31:0] = 32'd4294967295; 
    //             mask[95:64] = 32'd4294967295;   
    //             mult_ans = weight & mask; 
    //         end
    //         4'd6: begin
    //             mask = 128'b0;
    //             mask[95:32] = 32'd4294967295;   
    //             mult_ans = weight & mask; 
    //         end
    //         4'd7: begin
    //             mask = 128'b0;
    //             mask[95:0] = 64'd4294967295;   
    //             mult_ans = weight & mask; 
    //         end
    //         4'd8: begin
    //             mask = 128'b0;
    //             mask[127:96] = 32'd4294967295;   
    //             mult_ans = weight & mask; 
    //         end
    //         4'd9: begin
    //             mask = 128'b0;
    //             mask[127:96] = 32'd4294967295;  
    //             mask[31:0] = 32'd4294967295;
    //             mult_ans = weight & mask; 
    //         end
    //         4'd10: begin
    //             mask = 128'b0;
    //             mask[127:96] = 32'd4294967295;  
    //             mask[63:32] = 32'd4294967295;
    //             mult_ans = weight & mask; 
    //         end
    //         4'd11: begin
    //             mask = 128'b0;
    //             mask[127:96] = 32'd4294967295;  
    //             mask[63:0] = 64'd4294967295;
    //             mult_ans = weight & mask; 
    //         end
    //         4'd12: begin
    //             mask = 128'b0;
    //             mask[127:64] = 64'd4294967295;
    //             mult_ans = weight & mask; 
    //         end
    //         4'd13: begin
    //             mask = 128'b0;
    //             mask[127:96] = 32'd4294967295;  
    //             mask[31:0] = 32'd4294967295;
    //             mult_ans = weight & mask; 
    //         end
    //         4'd14: begin
    //             mask = 128'b0;
    //             mask[127:32] = 96'd4294967295;
    //             mult_ans = weight & mask; 
    //         end
    //         4'd15: begin
    //             mult_ans = weight;
    //         end
    //         default:    mult_ans = 4'bx;
    //     endcase
        
    //     // mult_output = mult_ans[31:0] + mult_ans[63:32] + mult_ans[95:64] + mult_ans[127:96];
    //     // mult_output = add_val3;
    // end

    // Addition_Subtraction add1(mult_ans[31:0], mult_ans[63:32], 1'b0, excpetion1, add_val1);
    // Addition_Subtraction add2(add_val1, mult_ans[95:64], 1'b0, excpetion2, add_val2);
    // Addition_Subtraction add3(add_val2, mult_ans[127:96], 1'b0, exception3, add_val3);

    // always@(add_val3 or spike_in) begin
    //     mult_output = add_val3;
    // end

endmodule