module (input wire [31:0] adder_potential, 
    input wire spiked, 
    output reg [31:0] potential_to_mem);

    // Reset if needed only, if not direct write

endmodule