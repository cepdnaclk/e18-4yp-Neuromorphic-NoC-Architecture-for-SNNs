module testbench_scaled;

    //neuron addresses
        source_addresses[129] = 12'd1024;        source_addresses[155] = 12'd1025;        source_addresses[156] = 12'd1026;        source_addresses[157] = 12'd1027;        source_addresses[158] = 12'd1028;        source_addresses[159] = 12'd1029;        source_addresses[182] = 12'd1030;        source_addresses[183] = 12'd1031;        source_addresses[184] = 12'd1032;        source_addresses[185] = 12'd1033;        source_addresses[186] = 12'd1034;        source_addresses[187] = 12'd1035;        source_addresses[209] = 12'd1036;        source_addresses[210] = 12'd1037;        source_addresses[211] = 12'd1038;        source_addresses[212] = 12'd1039;        source_addresses[213] = 12'd1040;        source_addresses[215] = 12'd1041;        source_addresses[216] = 12'd1042;        source_addresses[236] = 12'd1043;        source_addresses[237] = 12'd1044;        source_addresses[238] = 12'd1045;        source_addresses[239] = 12'd1046;        source_addresses[240] = 12'd1047;        source_addresses[241] = 12'd1048;        source_addresses[244] = 12'd1049;        source_addresses[263] = 12'd1050;        source_addresses[264] = 12'd1051;        source_addresses[265] = 12'd1052;        source_addresses[268] = 12'd1053;        source_addresses[269] = 12'd1054;        source_addresses[272] = 12'd1055;        source_addresses[290] = 12'd1056;        source_addresses[291] = 12'd1057;        source_addresses[292] = 12'd1058;        source_addresses[300] = 12'd1059;
        source_addresses[301] = 12'd1060;        source_addresses[318] = 12'd1061;        source_addresses[319] = 12'd1062;        source_addresses[320] = 12'd1063;        source_addresses[328] = 12'd1064;        source_addresses[329] = 12'd1065;        source_addresses[345] = 12'd1066;        source_addresses[346] = 12'd1067;        source_addresses[356] = 12'd1068;        source_addresses[357] = 12'd1069;        source_addresses[358] = 12'd1070;        source_addresses[372] = 12'd1071;        source_addresses[373] = 12'd1072;        source_addresses[384] = 12'd1073;        source_addresses[385] = 12'd1074;        source_addresses[386] = 12'd1075;        source_addresses[399] = 12'd1076;        source_addresses[400] = 12'd1077;
        source_addresses[412] = 12'd1078;        source_addresses[413] = 12'd1079;        source_addresses[414] = 12'd1080;        source_addresses[427] = 12'd1081;        source_addresses[428] = 12'd1082;        source_addresses[440] = 12'd1083;        source_addresses[441] = 12'd1084;        source_addresses[455] = 12'd1085;        source_addresses[456] = 12'd1086;        source_addresses[468] = 12'd1087;        source_addresses[483] = 12'd1088;        source_addresses[484] = 12'd1089;        source_addresses[495] = 12'd1090;        source_addresses[496] = 12'd1091;        source_addresses[511] = 12'd1092;        source_addresses[522] = 12'd1093;        source_addresses[539] = 12'd1094;        source_addresses[540] = 12'd1095;        source_addresses[548] = 12'd1096;        source_addresses[549] = 12'd1097;        source_addresses[567] = 12'd1098;        source_addresses[568] = 12'd1099;        source_addresses[574] = 12'd1100;        source_addresses[575] = 12'd1101;        source_addresses[576] = 12'd1102;        source_addresses[595] = 12'd1103;        source_addresses[596] = 12'd1104;        source_addresses[597] = 12'd1105;        source_addresses[598] = 12'd1106;        source_addresses[599] = 12'd1107;        source_addresses[600] = 12'd1108;
        source_addresses[601] = 12'd1109;        source_addresses[602] = 12'd1110;        source_addresses[603] = 12'd1111;        source_addresses[623] = 12'd1112;        source_addresses[624] = 12'd1113;        source_addresses[625] = 12'd1114;        source_addresses[626] = 12'd1115;        source_addresses[627] = 12'd1116;        source_addresses[628] = 12'd1117;        source_addresses[629] = 12'd1118;        source_addresses[653] = 12'd1119;        source_addresses[654] = 12'd1120;        source_addresses[655] = 12'd1121;