module network_interface_scaled (
        input wire spike0,
    input wire spike1,    input wire spike2,    input wire spike3,    input wire spike4,    input wire spike5,    input wire spike6,    input wire spike7,    input wire spike8,    input wire spike9,    input wire spike10,    input wire spike11,    input wire spike12,    input wire spike13,    input wire spike14,    input wire spike15,    input wire spike16,    input wire spike17,    input wire spike18,    input wire spike19,    input wire spike20,    input wire spike21,    input wire spike22,    input wire spike23,    input wire spike24,    input wire spike25,    input wire spike26,    input wire spike27,    input wire spike28,    input wire spike29,    input wire spike30,    input wire spike31,    input wire spike32,    input wire spike33,    input wire spike34,    input wire spike35,    input wire spike36,    input wire spike37,    input wire spike38,    input wire spike39,    input wire spike40,    input wire spike41,    input wire spike42,    input wire spike43,    input wire spike44,    input wire spike45,    input wire spike46,    input wire spike47,    input wire spike48,    input wire spike49,    input wire spike50,    input wire spike51,    input wire spike52,    input wire spike53,    input wire spike54,    input wire spike55,    input wire spike56,    input wire spike57,    input wire spike58,    input wire spike59,    input wire spike60,    input wire spike61,    input wire spike62,    input wire spike63,    input wire spike64,    input wire spike65,    input wire spike66,    input wire spike67,    input wire spike68,    input wire spike69,    input wire spike70,    input wire spike71,    input wire spike72,    input wire spike73,    input wire spike74,    input wire spike75,    input wire spike76,    input wire spike77,    input wire spike78,    input wire spike79,    input wire spike80,    input wire spike81,    input wire spike82,    input wire spike83,    input wire spike84,    input wire spike85,    input wire spike86,    input wire spike87,    input wire spike88,    input wire spike89,    input wire spike90,    input wire spike91,    input wire spike92,    input wire spike93,    input wire spike94,    input wire spike95,    input wire spike96,    input wire spike97,    input wire spike98,    input wire spike99,    input wire spike100,
    input wire spike101,    input wire spike102,    input wire spike103,    input wire spike104,    input wire spike105,    input wire spike106,    input wire spike107,    input wire spike108,    input wire spike109,    input wire spike110,    input wire spike111,    input wire spike112,    input wire spike113,    input wire spike114,    input wire spike115,    input wire spike116,    input wire spike117,    input wire spike118,    input wire spike119,    input wire spike120,    input wire spike121,    input wire spike122,    input wire spike123,    input wire spike124,    input wire spike125,    input wire spike126,    input wire spike127,    input wire spike128,    input wire spike129,    input wire spike130,    input wire spike131,    input wire spike132,    input wire spike133,    input wire spike134,    input wire spike135,    input wire spike136,    input wire spike137,    input wire spike138,    input wire spike139,    input wire spike140,    input wire spike141,    input wire spike142,    input wire spike143,    input wire spike144,    input wire spike145,    input wire spike146,    input wire spike147,    input wire spike148,    input wire spike149,    input wire spike150,    input wire spike151,    input wire spike152,    input wire spike153,    input wire spike154,    input wire spike155,    input wire spike156,    input wire spike157,    input wire spike158,    input wire spike159,    input wire spike160,    input wire spike161,    input wire spike162,    input wire spike163,    input wire spike164,    input wire spike165,    input wire spike166,    input wire spike167,    input wire spike168,    input wire spike169,    input wire spike170,    input wire spike171,    input wire spike172,    input wire spike173,    input wire spike174,    input wire spike175,    input wire spike176,    input wire spike177,    input wire spike178,    input wire spike179,    input wire spike180,    input wire spike181,    input wire spike182,    input wire spike183,    input wire spike184,    input wire spike185,    input wire spike186,    input wire spike187,    input wire spike188,    input wire spike189,    input wire spike190,    input wire spike191,    input wire spike192,    input wire spike193,    input wire spike194,    input wire spike195,    input wire spike196,    input wire spike197,    input wire spike198,    input wire spike199,    input wire spike200,
    input wire spike201,    input wire spike202,    input wire spike203,    input wire spike204,    input wire spike205,    input wire spike206,    input wire spike207,    input wire spike208,    input wire spike209,    input wire spike210,    input wire spike211,    input wire spike212,    input wire spike213,    input wire spike214,    input wire spike215,    input wire spike216,    input wire spike217,    input wire spike218,    input wire spike219,    input wire spike220,    input wire spike221,    input wire spike222,    input wire spike223,    input wire spike224,    input wire spike225,    input wire spike226,    input wire spike227,    input wire spike228,    input wire spike229,    input wire spike230,    input wire spike231,    input wire spike232,    input wire spike233,    input wire spike234,    input wire spike235,    input wire spike236,    input wire spike237,    input wire spike238,    input wire spike239,    input wire spike240,    input wire spike241,    input wire spike242,    input wire spike243,    input wire spike244,    input wire spike245,    input wire spike246,    input wire spike247,    input wire spike248,    input wire spike249,    input wire spike250,    input wire spike251,    input wire spike252,    input wire spike253,    input wire spike254,    input wire spike255,    input wire spike256,    input wire spike257,    input wire spike258,    input wire spike259,    input wire spike260,    input wire spike261,    input wire spike262,    input wire spike263,    input wire spike264,    input wire spike265,    input wire spike266,    input wire spike267,    input wire spike268,    input wire spike269,    input wire spike270,    input wire spike271,    input wire spike272,    input wire spike273,    input wire spike274,    input wire spike275,    input wire spike276,    input wire spike277,    input wire spike278,    input wire spike279,    input wire spike280,    input wire spike281,    input wire spike282,    input wire spike283,    input wire spike284,    input wire spike285,    input wire spike286,    input wire spike287,    input wire spike288,    input wire spike289,    input wire spike290,    input wire spike291,    input wire spike292,    input wire spike293,    input wire spike294,    input wire spike295,    input wire spike296,    input wire spike297,    input wire spike298,    input wire spike299,    input wire spike300,
    input wire spike301,    input wire spike302,    input wire spike303,    input wire spike304,    input wire spike305,    input wire spike306,    input wire spike307,    input wire spike308,    input wire spike309,    input wire spike310,    input wire spike311,    input wire spike312,    input wire spike313,    input wire spike314,    input wire spike315,    input wire spike316,    input wire spike317,    input wire spike318,    input wire spike319,    input wire spike320,    input wire spike321,    input wire spike322,    input wire spike323,    input wire spike324,    input wire spike325,    input wire spike326,    input wire spike327,    input wire spike328,    input wire spike329,    input wire spike330,    input wire spike331,    input wire spike332,    input wire spike333,    input wire spike334,    input wire spike335,    input wire spike336,    input wire spike337,    input wire spike338,    input wire spike339,    input wire spike340,    input wire spike341,    input wire spike342,    input wire spike343,    input wire spike344,    input wire spike345,    input wire spike346,    input wire spike347,    input wire spike348,    input wire spike349,    input wire spike350,    input wire spike351,    input wire spike352,    input wire spike353,    input wire spike354,    input wire spike355,    input wire spike356,    input wire spike357,    input wire spike358,    input wire spike359,    input wire spike360,    input wire spike361,    input wire spike362,    input wire spike363,    input wire spike364,    input wire spike365,    input wire spike366,    input wire spike367,    input wire spike368,    input wire spike369,    input wire spike370,    input wire spike371,    input wire spike372,    input wire spike373,    input wire spike374,    input wire spike375,    input wire spike376,    input wire spike377,    input wire spike378,    input wire spike379,    input wire spike380,    input wire spike381,    input wire spike382,    input wire spike383,    input wire spike384,    input wire spike385,    input wire spike386,    input wire spike387,    input wire spike388,    input wire spike389,    input wire spike390,    input wire spike391,    input wire spike392,    input wire spike393,    input wire spike394,    input wire spike395,    input wire spike396,    input wire spike397,    input wire spike398,    input wire spike399,    input wire spike400,
    input wire spike401,    input wire spike402,    input wire spike403,    input wire spike404,    input wire spike405,    input wire spike406,    input wire spike407,    input wire spike408,    input wire spike409,    input wire spike410,    input wire spike411,    input wire spike412,    input wire spike413,    input wire spike414,    input wire spike415,    input wire spike416,    input wire spike417,    input wire spike418,    input wire spike419,    input wire spike420,    input wire spike421,    input wire spike422,    input wire spike423,    input wire spike424,    input wire spike425,    input wire spike426,    input wire spike427,    input wire spike428,    input wire spike429,    input wire spike430,    input wire spike431,    input wire spike432,    input wire spike433,    input wire spike434,    input wire spike435,    input wire spike436,    input wire spike437,    input wire spike438,    input wire spike439,    input wire spike440,    input wire spike441,    input wire spike442,    input wire spike443,    input wire spike444,    input wire spike445,    input wire spike446,    input wire spike447,    input wire spike448,    input wire spike449,    input wire spike450,    input wire spike451,    input wire spike452,    input wire spike453,    input wire spike454,    input wire spike455,    input wire spike456,    input wire spike457,    input wire spike458,    input wire spike459,    input wire spike460,    input wire spike461,    input wire spike462,    input wire spike463,    input wire spike464,    input wire spike465,    input wire spike466,    input wire spike467,    input wire spike468,    input wire spike469,    input wire spike470,    input wire spike471,    input wire spike472,    input wire spike473,    input wire spike474,    input wire spike475,    input wire spike476,    input wire spike477,    input wire spike478,    input wire spike479,    input wire spike480,    input wire spike481,    input wire spike482,    input wire spike483,    input wire spike484,    input wire spike485,    input wire spike486,    input wire spike487,    input wire spike488,    input wire spike489,    input wire spike490,    input wire spike491,    input wire spike492,    input wire spike493,    input wire spike494,    input wire spike495,    input wire spike496,    input wire spike497,    input wire spike498,    input wire spike499,    input wire spike500,
    input wire spike501,    input wire spike502,    input wire spike503,    input wire spike504,    input wire spike505,    input wire spike506,    input wire spike507,    input wire spike508,    input wire spike509,    input wire spike510,    input wire spike511,    input wire spike512,    input wire spike513,    input wire spike514,    input wire spike515,    input wire spike516,    input wire spike517,    input wire spike518,    input wire spike519,    input wire spike520,    input wire spike521,    input wire spike522,    input wire spike523,    input wire spike524,    input wire spike525,    input wire spike526,    input wire spike527,    input wire spike528,    input wire spike529,    input wire spike530,    input wire spike531,    input wire spike532,    input wire spike533,    input wire spike534,    input wire spike535,    input wire spike536,    input wire spike537,    input wire spike538,    input wire spike539,    input wire spike540,    input wire spike541,    input wire spike542,    input wire spike543,    input wire spike544,    input wire spike545,    input wire spike546,    input wire spike547,    input wire spike548,    input wire spike549,    input wire spike550,    input wire spike551,    input wire spike552,    input wire spike553,    input wire spike554,    input wire spike555,    input wire spike556,    input wire spike557,    input wire spike558,    input wire spike559,    input wire spike560,    input wire spike561,    input wire spike562,    input wire spike563,    input wire spike564,    input wire spike565,    input wire spike566,    input wire spike567,    input wire spike568,    input wire spike569,    input wire spike570,    input wire spike571,    input wire spike572,    input wire spike573,    input wire spike574,    input wire spike575,    input wire spike576,    input wire spike577,    input wire spike578,    input wire spike579,    input wire spike580,    input wire spike581,    input wire spike582,    input wire spike583,    input wire spike584,    input wire spike585,    input wire spike586,    input wire spike587,    input wire spike588,    input wire spike589,    input wire spike590,    input wire spike591,    input wire spike592,    input wire spike593,    input wire spike594,    input wire spike595,    input wire spike596,    input wire spike597,    input wire spike598,    input wire spike599,    input wire spike600,
    input wire spike601,    input wire spike602,    input wire spike603,    input wire spike604,    input wire spike605,    input wire spike606,    input wire spike607,    input wire spike608,    input wire spike609,    input wire spike610,    input wire spike611,    input wire spike612,    input wire spike613,    input wire spike614,    input wire spike615,    input wire spike616,    input wire spike617,    input wire spike618,    input wire spike619,    input wire spike620,    input wire spike621,    input wire spike622,    input wire spike623,    input wire spike624,    input wire spike625,    input wire spike626,    input wire spike627,    input wire spike628,    input wire spike629,    input wire spike630,    input wire spike631,    input wire spike632,    input wire spike633,    input wire spike634,    input wire spike635,    input wire spike636,    input wire spike637,    input wire spike638,    input wire spike639,    input wire spike640,    input wire spike641,    input wire spike642,    input wire spike643,    input wire spike644,    input wire spike645,    input wire spike646,    input wire spike647,    input wire spike648,    input wire spike649,    input wire spike650,    input wire spike651,    input wire spike652,    input wire spike653,    input wire spike654,    input wire spike655,    input wire spike656,    input wire spike657,    input wire spike658,    input wire spike659,    input wire spike660,    input wire spike661,    input wire spike662,    input wire spike663,    input wire spike664,    input wire spike665,    input wire spike666,    input wire spike667,    input wire spike668,    input wire spike669,    input wire spike670,    input wire spike671,    input wire spike672,    input wire spike673,    input wire spike674,    input wire spike675,    input wire spike676,    input wire spike677,    input wire spike678,    input wire spike679,    input wire spike680,    input wire spike681,    input wire spike682,    input wire spike683,    input wire spike684,    input wire spike685,    input wire spike686,    input wire spike687,    input wire spike688,    input wire spike689,    input wire spike690,    input wire spike691,    input wire spike692,    input wire spike693,    input wire spike694,    input wire spike695,    input wire spike696,    input wire spike697,    input wire spike698,    input wire spike699,    input wire spike700,
    input wire spike701,    input wire spike702,    input wire spike703,    input wire spike704,    input wire spike705,    input wire spike706,    input wire spike707,    input wire spike708,    input wire spike709,    input wire spike710,    input wire spike711,    input wire spike712,    input wire spike713,    input wire spike714,    input wire spike715,    input wire spike716,    input wire spike717,    input wire spike718,    input wire spike719,    input wire spike720,    input wire spike721,    input wire spike722,    input wire spike723,    input wire spike724,    input wire spike725,    input wire spike726,    input wire spike727,    input wire spike728,    input wire spike729,    input wire spike730,    input wire spike731,    input wire spike732,    input wire spike733,    input wire spike734,    input wire spike735,    input wire spike736,    input wire spike737,    input wire spike738,    input wire spike739,    input wire spike740,    input wire spike741,    input wire spike742,    input wire spike743,    input wire spike744,    input wire spike745,    input wire spike746,    input wire spike747,    input wire spike748,    input wire spike749,    input wire spike750,    input wire spike751,    input wire spike752,    input wire spike753,    input wire spike754,    input wire spike755,    input wire spike756,    input wire spike757,    input wire spike758,    input wire spike759,    input wire spike760,    input wire spike761,    input wire spike762,    input wire spike763,    input wire spike764,    input wire spike765,    input wire spike766,    input wire spike767,    input wire spike768,    input wire spike769,    input wire spike770,    input wire spike771,    input wire spike772,    input wire spike773,    input wire spike774,    input wire spike775,    input wire spike776,    input wire spike777,    input wire spike778,    input wire spike779,    input wire spike780,    input wire spike781,    input wire spike782,    input wire spike783,    input wire spike784,    input wire spike785,    input wire spike786,    input wire spike787,    input wire spike788,    input wire spike789,    input wire spike790,    input wire spike791,    input wire spike792,    input wire spike793,    input wire spike794,    input wire spike795,    input wire spike796,    input wire spike797,    input wire spike798,    input wire spike799,    input wire spike800,
    input wire spike801,    input wire spike802,    input wire spike803,    input wire spike804,    input wire spike805,    input wire spike806,    input wire spike807,    input wire spike808,    input wire spike809,    input wire spike810,    input wire spike811,    input wire spike812,    input wire spike813,    input wire spike814,    input wire spike815,    input wire spike816,    input wire spike817,    input wire spike818,    input wire spike819,    input wire spike820,    input wire spike821,    input wire spike822,    input wire spike823,    input wire spike824,    input wire spike825,    input wire spike826,    input wire spike827,    input wire spike828,    input wire spike829,    input wire spike830,    input wire spike831,    input wire spike832,    input wire spike833,    input wire spike834,    input wire spike835,    input wire spike836,    input wire spike837,    input wire spike838,    input wire spike839,    input wire spike840,    input wire spike841,    input wire spike842,    input wire spike843,    input wire spike844,    input wire spike845,    input wire spike846,    input wire spike847,    input wire spike848,    input wire spike849,    input wire spike850,    input wire spike851,    input wire spike852,    input wire spike853,    input wire spike854,    input wire spike855,    input wire spike856,    input wire spike857,    input wire spike858,    input wire spike859,    input wire spike860,    input wire spike861,    input wire spike862,    input wire spike863,    input wire spike864,    input wire spike865,    input wire spike866,    input wire spike867,    input wire spike868,    input wire spike869,    input wire spike870,    input wire spike871,    input wire spike872,    input wire spike873,    input wire spike874,    input wire spike875,    input wire spike876,    input wire spike877,    input wire spike878,    input wire spike879,    input wire spike880,    input wire spike881,    input wire spike882,    input wire spike883,    input wire spike884,    input wire spike885,    input wire spike886,    input wire spike887,    input wire spike888,    input wire spike889,    input wire spike890,    input wire spike891,    input wire spike892,    input wire spike893,    input wire spike894,    input wire spike895,    input wire spike896,    input wire spike897,    input wire spike898,    input wire spike899,    input wire spike900,
    input wire spike901,    input wire spike902,    input wire spike903,    input wire spike904,    input wire spike905,    input wire spike906,    input wire spike907,    input wire spike908,    input wire spike909,    input wire spike910,    input wire spike911,    input wire spike912,    input wire spike913,    input wire spike914,    input wire spike915,    input wire spike916,    input wire spike917,    input wire spike918,    input wire spike919,    input wire spike920,    input wire spike921,    input wire spike922,    input wire spike923,    input wire spike924,    input wire spike925,    input wire spike926,    input wire spike927,    input wire spike928,    input wire spike929,    input wire spike930,    input wire spike931,    input wire spike932,    input wire spike933,    input wire spike934,    input wire spike935,    input wire spike936,    input wire spike937,    input wire spike938,    input wire spike939,    input wire spike940,    input wire spike941,    input wire spike942,    input wire spike943,    input wire spike944,    input wire spike945,    input wire spike946,    input wire spike947,    input wire spike948,    input wire spike949,    input wire spike950,    input wire spike951,    input wire spike952,    input wire spike953,    input wire spike954,    input wire spike955,    input wire spike956,    input wire spike957,    input wire spike958,    input wire spike959,    input wire spike960,    input wire spike961,    input wire spike962,    input wire spike963,    input wire spike964,    input wire spike965,    input wire spike966,    input wire spike967,    input wire spike968,    input wire spike969,    input wire spike970,    input wire spike971,    input wire spike972,    input wire spike973,    input wire spike974,    input wire spike975,    input wire spike976,    input wire spike977,    input wire spike978,    input wire spike979,    input wire spike980,    input wire spike981,    input wire spike982,    input wire spike983,    input wire spike984,    input wire spike985,    input wire spike986,    input wire spike987,    input wire spike988,    input wire spike989,    input wire spike990,    input wire spike991,    input wire spike992,    input wire spike993,    input wire spike994,    input wire spike995,    input wire spike996,    input wire spike997,    input wire spike998,    input wire spike999,    input wire spike1000,
    input wire spike1001,    input wire spike1002,    input wire spike1003,    input wire spike1004,    input wire spike1005,    input wire spike1006,    input wire spike1007,    input wire spike1008,    input wire spike1009,    input wire spike1010,    input wire spike1011,    input wire spike1012,    input wire spike1013,    input wire spike1014,    input wire spike1015,    input wire spike1016,    input wire spike1017,    input wire spike1018,    input wire spike1019,    input wire spike1020,    input wire spike1021,    input wire spike1022,    input wire spike1023,
output reg[11:0]     spike_out_source0,
    spike_out_source1,    spike_out_source2,    spike_out_source3,    spike_out_source4,    spike_out_source5,    spike_out_source6,    spike_out_source7,    spike_out_source8,    spike_out_source9,    spike_out_source10,    spike_out_source11,    spike_out_source12,    spike_out_source13,    spike_out_source14,    spike_out_source15,    spike_out_source16,    spike_out_source17,    spike_out_source18,    spike_out_source19,    spike_out_source20,    spike_out_source21,    spike_out_source22,    spike_out_source23,    spike_out_source24,    spike_out_source25,    spike_out_source26,    spike_out_source27,    spike_out_source28,    spike_out_source29,    spike_out_source30,    spike_out_source31,    spike_out_source32,    spike_out_source33,    spike_out_source34,    spike_out_source35,    spike_out_source36,    spike_out_source37,    spike_out_source38,    spike_out_source39,    spike_out_source40,    spike_out_source41,    spike_out_source42,    spike_out_source43,    spike_out_source44,    spike_out_source45,    spike_out_source46,    spike_out_source47,    spike_out_source48,    spike_out_source49,    spike_out_source50,    spike_out_source51,    spike_out_source52,    spike_out_source53,    spike_out_source54,    spike_out_source55,    spike_out_source56,    spike_out_source57,    spike_out_source58,    spike_out_source59,    spike_out_source60,    spike_out_source61,    spike_out_source62,    spike_out_source63,    spike_out_source64,    spike_out_source65,    spike_out_source66,    spike_out_source67,    spike_out_source68,    spike_out_source69,    spike_out_source70,    spike_out_source71,    spike_out_source72,    spike_out_source73,    spike_out_source74,    spike_out_source75,    spike_out_source76,    spike_out_source77,    spike_out_source78,    spike_out_source79,    spike_out_source80,    spike_out_source81,    spike_out_source82,    spike_out_source83,    spike_out_source84,    spike_out_source85,    spike_out_source86,    spike_out_source87,    spike_out_source88,    spike_out_source89,    spike_out_source90,    spike_out_source91,    spike_out_source92,    spike_out_source93,    spike_out_source94,    spike_out_source95,    spike_out_source96,    spike_out_source97,    spike_out_source98,    spike_out_source99,    spike_out_source100,
    spike_out_source101,    spike_out_source102,    spike_out_source103,    spike_out_source104,    spike_out_source105,    spike_out_source106,    spike_out_source107,    spike_out_source108,    spike_out_source109,    spike_out_source110,    spike_out_source111,    spike_out_source112,    spike_out_source113,    spike_out_source114,    spike_out_source115,    spike_out_source116,    spike_out_source117,    spike_out_source118,    spike_out_source119,    spike_out_source120,    spike_out_source121,    spike_out_source122,    spike_out_source123,    spike_out_source124,    spike_out_source125,    spike_out_source126,    spike_out_source127,    spike_out_source128,    spike_out_source129,    spike_out_source130,    spike_out_source131,    spike_out_source132,    spike_out_source133,    spike_out_source134,    spike_out_source135,    spike_out_source136,    spike_out_source137,    spike_out_source138,    spike_out_source139,    spike_out_source140,    spike_out_source141,    spike_out_source142,    spike_out_source143,    spike_out_source144,    spike_out_source145,    spike_out_source146,    spike_out_source147,    spike_out_source148,    spike_out_source149,    spike_out_source150,    spike_out_source151,    spike_out_source152,    spike_out_source153,    spike_out_source154,    spike_out_source155,    spike_out_source156,    spike_out_source157,    spike_out_source158,    spike_out_source159,    spike_out_source160,    spike_out_source161,    spike_out_source162,    spike_out_source163,    spike_out_source164,    spike_out_source165,    spike_out_source166,    spike_out_source167,    spike_out_source168,    spike_out_source169,    spike_out_source170,    spike_out_source171,    spike_out_source172,    spike_out_source173,    spike_out_source174,    spike_out_source175,    spike_out_source176,    spike_out_source177,    spike_out_source178,    spike_out_source179,    spike_out_source180,    spike_out_source181,    spike_out_source182,    spike_out_source183,    spike_out_source184,    spike_out_source185,    spike_out_source186,    spike_out_source187,    spike_out_source188,    spike_out_source189,    spike_out_source190,    spike_out_source191,    spike_out_source192,    spike_out_source193,    spike_out_source194,    spike_out_source195,    spike_out_source196,    spike_out_source197,    spike_out_source198,    spike_out_source199,    spike_out_source200,
    spike_out_source201,    spike_out_source202,    spike_out_source203,    spike_out_source204,    spike_out_source205,    spike_out_source206,    spike_out_source207,    spike_out_source208,    spike_out_source209,    spike_out_source210,    spike_out_source211,    spike_out_source212,    spike_out_source213,    spike_out_source214,    spike_out_source215,    spike_out_source216,    spike_out_source217,    spike_out_source218,    spike_out_source219,    spike_out_source220,    spike_out_source221,    spike_out_source222,    spike_out_source223,    spike_out_source224,    spike_out_source225,    spike_out_source226,    spike_out_source227,    spike_out_source228,    spike_out_source229,    spike_out_source230,    spike_out_source231,    spike_out_source232,    spike_out_source233,    spike_out_source234,    spike_out_source235,    spike_out_source236,    spike_out_source237,    spike_out_source238,    spike_out_source239,    spike_out_source240,    spike_out_source241,    spike_out_source242,    spike_out_source243,    spike_out_source244,    spike_out_source245,    spike_out_source246,    spike_out_source247,    spike_out_source248,    spike_out_source249,    spike_out_source250,    spike_out_source251,    spike_out_source252,    spike_out_source253,    spike_out_source254,    spike_out_source255,    spike_out_source256,    spike_out_source257,    spike_out_source258,    spike_out_source259,    spike_out_source260,    spike_out_source261,    spike_out_source262,    spike_out_source263,    spike_out_source264,    spike_out_source265,    spike_out_source266,    spike_out_source267,    spike_out_source268,    spike_out_source269,    spike_out_source270,    spike_out_source271,    spike_out_source272,    spike_out_source273,    spike_out_source274,    spike_out_source275,    spike_out_source276,    spike_out_source277,    spike_out_source278,    spike_out_source279,    spike_out_source280,    spike_out_source281,    spike_out_source282,    spike_out_source283,    spike_out_source284,    spike_out_source285,    spike_out_source286,    spike_out_source287,    spike_out_source288,    spike_out_source289,    spike_out_source290,    spike_out_source291,    spike_out_source292,    spike_out_source293,    spike_out_source294,    spike_out_source295,    spike_out_source296,    spike_out_source297,    spike_out_source298,    spike_out_source299,    spike_out_source300,
    spike_out_source301,    spike_out_source302,    spike_out_source303,    spike_out_source304,    spike_out_source305,    spike_out_source306,    spike_out_source307,    spike_out_source308,    spike_out_source309,    spike_out_source310,    spike_out_source311,    spike_out_source312,    spike_out_source313,    spike_out_source314,    spike_out_source315,    spike_out_source316,    spike_out_source317,    spike_out_source318,    spike_out_source319,    spike_out_source320,    spike_out_source321,    spike_out_source322,    spike_out_source323,    spike_out_source324,    spike_out_source325,    spike_out_source326,    spike_out_source327,    spike_out_source328,    spike_out_source329,    spike_out_source330,    spike_out_source331,    spike_out_source332,    spike_out_source333,    spike_out_source334,    spike_out_source335,    spike_out_source336,    spike_out_source337,    spike_out_source338,    spike_out_source339,    spike_out_source340,    spike_out_source341,    spike_out_source342,    spike_out_source343,    spike_out_source344,    spike_out_source345,    spike_out_source346,    spike_out_source347,    spike_out_source348,    spike_out_source349,    spike_out_source350,    spike_out_source351,    spike_out_source352,    spike_out_source353,    spike_out_source354,    spike_out_source355,    spike_out_source356,    spike_out_source357,    spike_out_source358,    spike_out_source359,    spike_out_source360,    spike_out_source361,    spike_out_source362,    spike_out_source363,    spike_out_source364,    spike_out_source365,    spike_out_source366,    spike_out_source367,    spike_out_source368,    spike_out_source369,    spike_out_source370,    spike_out_source371,    spike_out_source372,    spike_out_source373,    spike_out_source374,    spike_out_source375,    spike_out_source376,    spike_out_source377,    spike_out_source378,    spike_out_source379,    spike_out_source380,    spike_out_source381,    spike_out_source382,    spike_out_source383,    spike_out_source384,    spike_out_source385,    spike_out_source386,    spike_out_source387,    spike_out_source388,    spike_out_source389,    spike_out_source390,    spike_out_source391,    spike_out_source392,    spike_out_source393,    spike_out_source394,    spike_out_source395,    spike_out_source396,    spike_out_source397,    spike_out_source398,    spike_out_source399,    spike_out_source400,
    spike_out_source401,    spike_out_source402,    spike_out_source403,    spike_out_source404,    spike_out_source405,    spike_out_source406,    spike_out_source407,    spike_out_source408,    spike_out_source409,    spike_out_source410,    spike_out_source411,    spike_out_source412,    spike_out_source413,    spike_out_source414,    spike_out_source415,    spike_out_source416,    spike_out_source417,    spike_out_source418,    spike_out_source419,    spike_out_source420,    spike_out_source421,    spike_out_source422,    spike_out_source423,    spike_out_source424,    spike_out_source425,    spike_out_source426,    spike_out_source427,    spike_out_source428,    spike_out_source429,    spike_out_source430,    spike_out_source431,    spike_out_source432,    spike_out_source433,    spike_out_source434,    spike_out_source435,    spike_out_source436,    spike_out_source437,    spike_out_source438,    spike_out_source439,    spike_out_source440,    spike_out_source441,    spike_out_source442,    spike_out_source443,    spike_out_source444,    spike_out_source445,    spike_out_source446,    spike_out_source447,    spike_out_source448,    spike_out_source449,    spike_out_source450,    spike_out_source451,    spike_out_source452,    spike_out_source453,    spike_out_source454,    spike_out_source455,    spike_out_source456,    spike_out_source457,    spike_out_source458,    spike_out_source459,    spike_out_source460,    spike_out_source461,    spike_out_source462,    spike_out_source463,    spike_out_source464,    spike_out_source465,    spike_out_source466,    spike_out_source467,    spike_out_source468,    spike_out_source469,    spike_out_source470,    spike_out_source471,    spike_out_source472,    spike_out_source473,    spike_out_source474,    spike_out_source475,    spike_out_source476,    spike_out_source477,    spike_out_source478,    spike_out_source479,    spike_out_source480,    spike_out_source481,    spike_out_source482,    spike_out_source483,    spike_out_source484,    spike_out_source485,    spike_out_source486,    spike_out_source487,    spike_out_source488,    spike_out_source489,    spike_out_source490,    spike_out_source491,    spike_out_source492,    spike_out_source493,    spike_out_source494,    spike_out_source495,    spike_out_source496,    spike_out_source497,    spike_out_source498,    spike_out_source499,    spike_out_source500,
    spike_out_source501,    spike_out_source502,    spike_out_source503,    spike_out_source504,    spike_out_source505,    spike_out_source506,    spike_out_source507,    spike_out_source508,    spike_out_source509,    spike_out_source510,    spike_out_source511,    spike_out_source512,    spike_out_source513,    spike_out_source514,    spike_out_source515,    spike_out_source516,    spike_out_source517,    spike_out_source518,    spike_out_source519,    spike_out_source520,    spike_out_source521,    spike_out_source522,    spike_out_source523,    spike_out_source524,    spike_out_source525,    spike_out_source526,    spike_out_source527,    spike_out_source528,    spike_out_source529,    spike_out_source530,    spike_out_source531,    spike_out_source532,    spike_out_source533,    spike_out_source534,    spike_out_source535,    spike_out_source536,    spike_out_source537,    spike_out_source538,    spike_out_source539,    spike_out_source540,    spike_out_source541,    spike_out_source542,    spike_out_source543,    spike_out_source544,    spike_out_source545,    spike_out_source546,    spike_out_source547,    spike_out_source548,    spike_out_source549,    spike_out_source550,    spike_out_source551,    spike_out_source552,    spike_out_source553,    spike_out_source554,    spike_out_source555,    spike_out_source556,    spike_out_source557,    spike_out_source558,    spike_out_source559,    spike_out_source560,    spike_out_source561,    spike_out_source562,    spike_out_source563,    spike_out_source564,    spike_out_source565,    spike_out_source566,    spike_out_source567,    spike_out_source568,    spike_out_source569,    spike_out_source570,    spike_out_source571,    spike_out_source572,    spike_out_source573,    spike_out_source574,    spike_out_source575,    spike_out_source576,    spike_out_source577,    spike_out_source578,    spike_out_source579,    spike_out_source580,    spike_out_source581,    spike_out_source582,    spike_out_source583,    spike_out_source584,    spike_out_source585,    spike_out_source586,    spike_out_source587,    spike_out_source588,    spike_out_source589,    spike_out_source590,    spike_out_source591,    spike_out_source592,    spike_out_source593,    spike_out_source594,    spike_out_source595,    spike_out_source596,    spike_out_source597,    spike_out_source598,    spike_out_source599,    spike_out_source600,
    spike_out_source601,    spike_out_source602,    spike_out_source603,    spike_out_source604,    spike_out_source605,    spike_out_source606,    spike_out_source607,    spike_out_source608,    spike_out_source609,    spike_out_source610,    spike_out_source611,    spike_out_source612,    spike_out_source613,    spike_out_source614,    spike_out_source615,    spike_out_source616,    spike_out_source617,    spike_out_source618,    spike_out_source619,    spike_out_source620,    spike_out_source621,    spike_out_source622,    spike_out_source623,    spike_out_source624,    spike_out_source625,    spike_out_source626,    spike_out_source627,    spike_out_source628,    spike_out_source629,    spike_out_source630,    spike_out_source631,    spike_out_source632,    spike_out_source633,    spike_out_source634,    spike_out_source635,    spike_out_source636,    spike_out_source637,    spike_out_source638,    spike_out_source639,    spike_out_source640,    spike_out_source641,    spike_out_source642,    spike_out_source643,    spike_out_source644,    spike_out_source645,    spike_out_source646,    spike_out_source647,    spike_out_source648,    spike_out_source649,    spike_out_source650,    spike_out_source651,    spike_out_source652,    spike_out_source653,    spike_out_source654,    spike_out_source655,    spike_out_source656,    spike_out_source657,    spike_out_source658,    spike_out_source659,    spike_out_source660,    spike_out_source661,    spike_out_source662,    spike_out_source663,    spike_out_source664,    spike_out_source665,    spike_out_source666,    spike_out_source667,    spike_out_source668,    spike_out_source669,    spike_out_source670,    spike_out_source671,    spike_out_source672,    spike_out_source673,    spike_out_source674,    spike_out_source675,    spike_out_source676,    spike_out_source677,    spike_out_source678,    spike_out_source679,    spike_out_source680,    spike_out_source681,    spike_out_source682,    spike_out_source683,    spike_out_source684,    spike_out_source685,    spike_out_source686,    spike_out_source687,    spike_out_source688,    spike_out_source689,    spike_out_source690,    spike_out_source691,    spike_out_source692,    spike_out_source693,    spike_out_source694,    spike_out_source695,    spike_out_source696,    spike_out_source697,    spike_out_source698,    spike_out_source699,    spike_out_source700,
    spike_out_source701,    spike_out_source702,    spike_out_source703,    spike_out_source704,    spike_out_source705,    spike_out_source706,    spike_out_source707,    spike_out_source708,    spike_out_source709,    spike_out_source710,    spike_out_source711,    spike_out_source712,    spike_out_source713,    spike_out_source714,    spike_out_source715,    spike_out_source716,    spike_out_source717,    spike_out_source718,    spike_out_source719,    spike_out_source720,    spike_out_source721,    spike_out_source722,    spike_out_source723,    spike_out_source724,    spike_out_source725,    spike_out_source726,    spike_out_source727,    spike_out_source728,    spike_out_source729,    spike_out_source730,    spike_out_source731,    spike_out_source732,    spike_out_source733,    spike_out_source734,    spike_out_source735,    spike_out_source736,    spike_out_source737,    spike_out_source738,    spike_out_source739,    spike_out_source740,    spike_out_source741,    spike_out_source742,    spike_out_source743,    spike_out_source744,    spike_out_source745,    spike_out_source746,    spike_out_source747,    spike_out_source748,    spike_out_source749,    spike_out_source750,    spike_out_source751,    spike_out_source752,    spike_out_source753,    spike_out_source754,    spike_out_source755,    spike_out_source756,    spike_out_source757,    spike_out_source758,    spike_out_source759,    spike_out_source760,    spike_out_source761,    spike_out_source762,    spike_out_source763,    spike_out_source764,    spike_out_source765,    spike_out_source766,    spike_out_source767,    spike_out_source768,    spike_out_source769,    spike_out_source770,    spike_out_source771,    spike_out_source772,    spike_out_source773,    spike_out_source774,    spike_out_source775,    spike_out_source776,    spike_out_source777,    spike_out_source778,    spike_out_source779,    spike_out_source780,    spike_out_source781,    spike_out_source782,    spike_out_source783,    spike_out_source784,    spike_out_source785,    spike_out_source786,    spike_out_source787,    spike_out_source788,    spike_out_source789,    spike_out_source790,    spike_out_source791,    spike_out_source792,    spike_out_source793,    spike_out_source794,    spike_out_source795,    spike_out_source796,    spike_out_source797,    spike_out_source798,    spike_out_source799,    spike_out_source800,
    spike_out_source801,    spike_out_source802,    spike_out_source803,    spike_out_source804,    spike_out_source805,    spike_out_source806,    spike_out_source807,    spike_out_source808,    spike_out_source809,    spike_out_source810,    spike_out_source811,    spike_out_source812,    spike_out_source813,    spike_out_source814,    spike_out_source815,    spike_out_source816,    spike_out_source817,    spike_out_source818,    spike_out_source819,    spike_out_source820,    spike_out_source821,    spike_out_source822,    spike_out_source823,    spike_out_source824,    spike_out_source825,    spike_out_source826,    spike_out_source827,    spike_out_source828,    spike_out_source829,    spike_out_source830,    spike_out_source831,    spike_out_source832,    spike_out_source833,    spike_out_source834,    spike_out_source835,    spike_out_source836,    spike_out_source837,    spike_out_source838,    spike_out_source839,    spike_out_source840,    spike_out_source841,    spike_out_source842,    spike_out_source843,    spike_out_source844,    spike_out_source845,    spike_out_source846,    spike_out_source847,    spike_out_source848,    spike_out_source849,    spike_out_source850,    spike_out_source851,    spike_out_source852,    spike_out_source853,    spike_out_source854,    spike_out_source855,    spike_out_source856,    spike_out_source857,    spike_out_source858,    spike_out_source859,    spike_out_source860,    spike_out_source861,    spike_out_source862,    spike_out_source863,    spike_out_source864,    spike_out_source865,    spike_out_source866,    spike_out_source867,    spike_out_source868,    spike_out_source869,    spike_out_source870,    spike_out_source871,    spike_out_source872,    spike_out_source873,    spike_out_source874,    spike_out_source875,    spike_out_source876,    spike_out_source877,    spike_out_source878,    spike_out_source879,    spike_out_source880,    spike_out_source881,    spike_out_source882,    spike_out_source883,    spike_out_source884,    spike_out_source885,    spike_out_source886,    spike_out_source887,    spike_out_source888,    spike_out_source889,    spike_out_source890,    spike_out_source891,    spike_out_source892,    spike_out_source893,    spike_out_source894,    spike_out_source895,    spike_out_source896,    spike_out_source897,    spike_out_source898,    spike_out_source899,    spike_out_source900,
    spike_out_source901,    spike_out_source902,    spike_out_source903,    spike_out_source904,    spike_out_source905,    spike_out_source906,    spike_out_source907,    spike_out_source908,    spike_out_source909,    spike_out_source910,    spike_out_source911,    spike_out_source912,    spike_out_source913,    spike_out_source914,    spike_out_source915,    spike_out_source916,    spike_out_source917,    spike_out_source918,    spike_out_source919,    spike_out_source920,    spike_out_source921,    spike_out_source922,    spike_out_source923,    spike_out_source924,    spike_out_source925,    spike_out_source926,    spike_out_source927,    spike_out_source928,    spike_out_source929,    spike_out_source930,    spike_out_source931,    spike_out_source932,    spike_out_source933,    spike_out_source934,    spike_out_source935,    spike_out_source936,    spike_out_source937,    spike_out_source938,    spike_out_source939,    spike_out_source940,    spike_out_source941,    spike_out_source942,    spike_out_source943,    spike_out_source944,    spike_out_source945,    spike_out_source946,    spike_out_source947,    spike_out_source948,    spike_out_source949,    spike_out_source950,    spike_out_source951,    spike_out_source952,    spike_out_source953,    spike_out_source954,    spike_out_source955,    spike_out_source956,    spike_out_source957,    spike_out_source958,    spike_out_source959,    spike_out_source960,    spike_out_source961,    spike_out_source962,    spike_out_source963,    spike_out_source964,    spike_out_source965,    spike_out_source966,    spike_out_source967,    spike_out_source968,    spike_out_source969,    spike_out_source970,    spike_out_source971,    spike_out_source972,    spike_out_source973,    spike_out_source974,    spike_out_source975,    spike_out_source976,    spike_out_source977,    spike_out_source978,    spike_out_source979,    spike_out_source980,    spike_out_source981,    spike_out_source982,    spike_out_source983,    spike_out_source984,    spike_out_source985,    spike_out_source986,    spike_out_source987,    spike_out_source988,    spike_out_source989,    spike_out_source990,    spike_out_source991,    spike_out_source992,    spike_out_source993,    spike_out_source994,    spike_out_source995,    spike_out_source996,    spike_out_source997,    spike_out_source998,    spike_out_source999,    spike_out_source1000,
    spike_out_source1001,    spike_out_source1002,    spike_out_source1003,    spike_out_source1004,    spike_out_source1005,    spike_out_source1006,    spike_out_source1007,    spike_out_source1008,    spike_out_source1009,    spike_out_source1010,    spike_out_source1011,    spike_out_source1012,    spike_out_source1013,    spike_out_source1014,    spike_out_source1015,    spike_out_source1016,    spike_out_source1017,    spike_out_source1018,    spike_out_source1019,    spike_out_source1020,    spike_out_source1021,    spike_out_source1022,    spike_out_source1023,
    output wire output
);

    parameter number_of_neurons= 1024;
    reg spike_register[0:number_of_neurons-1];
    always @(clear, lock1, spike0, spike1, spike2, spike3, spike4, spike5, spike6, spike7, spike8, spike9, spike10, spike11, spike12, spike13, spike14, spike15, spike16, spike17, spike18, spike19, spike20, spike21, spike22, spike23, spike24, spike25, spike26, spike27, spike28, spike29, spike30, spike31, spike32, spike33, spike34, spike35, spike36, spike37, spike38, spike39, spike40, spike41, spike42, spike43, spike44, spike45, spike46, spike47, spike48, spike49) begin
        spike_register[0] = spike0;

        spike_register[1] = spike1;        spike_register[2] = spike2;        spike_register[3] = spike3;        spike_register[4] = spike4;        spike_register[5] = spike5;        spike_register[6] = spike6;        spike_register[7] = spike7;        spike_register[8] = spike8;        spike_register[9] = spike9;        spike_register[10] = spike10;        spike_register[11] = spike11;        spike_register[12] = spike12;        spike_register[13] = spike13;        spike_register[14] = spike14;        spike_register[15] = spike15;        spike_register[16] = spike16;        spike_register[17] = spike17;        spike_register[18] = spike18;        spike_register[19] = spike19;        spike_register[20] = spike20;        spike_register[21] = spike21;        spike_register[22] = spike22;        spike_register[23] = spike23;        spike_register[24] = spike24;        spike_register[25] = spike25;        spike_register[26] = spike26;        spike_register[27] = spike27;        spike_register[28] = spike28;        spike_register[29] = spike29;        spike_register[30] = spike30;        spike_register[31] = spike31;        spike_register[32] = spike32;        spike_register[33] = spike33;        spike_register[34] = spike34;        spike_register[35] = spike35;        spike_register[36] = spike36;        spike_register[37] = spike37;        spike_register[38] = spike38;        spike_register[39] = spike39;        spike_register[40] = spike40;        spike_register[41] = spike41;        spike_register[42] = spike42;        spike_register[43] = spike43;        spike_register[44] = spike44;        spike_register[45] = spike45;        spike_register[46] = spike46;        spike_register[47] = spike47;        spike_register[48] = spike48;        spike_register[49] = spike49;
        #0.5
        if(clear == 1'b0) begin
            for(i1 = 0; i1 <=49; i1= i1+1) begin
                if(spike_register[i1] == 1 && lock1 == 0) begin
                    lock1 = 1;
                    for(j1 = connection_pointer[i1]; j1 < connection_pointer[i1+1]; j1= j1+1) begin
                        packet1 = #0.1 {neuron_addresses[i1], downstream_connections[j1]};
                    end
                    spike_register[i1] = 0;
                    lock1 = 0;
                end
            end
        end

    end
    always @(clear, lock2, spike50, spike51, spike52, spike53, spike54, spike55, spike56, spike57, spike58, spike59, spike60, spike61, spike62, spike63, spike64, spike65, spike66, spike67, spike68, spike69, spike70, spike71, spike72, spike73, spike74, spike75, spike76, spike77, spike78, spike79, spike80, spike81, spike82, spike83, spike84, spike85, spike86, spike87, spike88, spike89, spike90, spike91, spike92, spike93, spike94, spike95, spike96, spike97, spike98, spike99) begin
        spike_register[50] = spike50;        spike_register[51] = spike51;        spike_register[52] = spike52;        spike_register[53] = spike53;        spike_register[54] = spike54;        spike_register[55] = spike55;        spike_register[56] = spike56;        spike_register[57] = spike57;        spike_register[58] = spike58;        spike_register[59] = spike59;        spike_register[60] = spike60;        spike_register[61] = spike61;        spike_register[62] = spike62;        spike_register[63] = spike63;        spike_register[64] = spike64;        spike_register[65] = spike65;        spike_register[66] = spike66;        spike_register[67] = spike67;        spike_register[68] = spike68;        spike_register[69] = spike69;        spike_register[70] = spike70;        spike_register[71] = spike71;        spike_register[72] = spike72;        spike_register[73] = spike73;        spike_register[74] = spike74;        spike_register[75] = spike75;        spike_register[76] = spike76;        spike_register[77] = spike77;        spike_register[78] = spike78;        spike_register[79] = spike79;        spike_register[80] = spike80;        spike_register[81] = spike81;        spike_register[82] = spike82;        spike_register[83] = spike83;        spike_register[84] = spike84;        spike_register[85] = spike85;        spike_register[86] = spike86;        spike_register[87] = spike87;        spike_register[88] = spike88;        spike_register[89] = spike89;        spike_register[90] = spike90;        spike_register[91] = spike91;        spike_register[92] = spike92;        spike_register[93] = spike93;        spike_register[94] = spike94;        spike_register[95] = spike95;        spike_register[96] = spike96;        spike_register[97] = spike97;        spike_register[98] = spike98;        spike_register[99] = spike99;
        #0.5
        if(clear == 1'b0) begin
            for(i2 = 50; i2 <=99; i2= i2+1) begin
                if(spike_register[i2] == 1 && lock2 == 0) begin
                    lock2 = 1;
                    for(j2 = connection_pointer[i2]; j2 < connection_pointer[i2+1]; j2= j2+1) begin
                        packet2 = #0.1 {neuron_addresses[i2], downstream_connections[j2]};
                    end
                    spike_register[i2] = 0;
                    lock2 = 0;
                end
            end
        end

    end
    always @(clear, lock3, spike100, spike101, spike102, spike103, spike104, spike105, spike106, spike107, spike108, spike109, spike110, spike111, spike112, spike113, spike114, spike115, spike116, spike117, spike118, spike119, spike120, spike121, spike122, spike123, spike124, spike125, spike126, spike127, spike128, spike129, spike130, spike131, spike132, spike133, spike134, spike135, spike136, spike137, spike138, spike139, spike140, spike141, spike142, spike143, spike144, spike145, spike146, spike147, spike148, spike149) begin
        spike_register[100] = spike100;

        spike_register[101] = spike101;        spike_register[102] = spike102;        spike_register[103] = spike103;        spike_register[104] = spike104;        spike_register[105] = spike105;        spike_register[106] = spike106;        spike_register[107] = spike107;        spike_register[108] = spike108;        spike_register[109] = spike109;        spike_register[110] = spike110;        spike_register[111] = spike111;        spike_register[112] = spike112;        spike_register[113] = spike113;        spike_register[114] = spike114;        spike_register[115] = spike115;        spike_register[116] = spike116;        spike_register[117] = spike117;        spike_register[118] = spike118;        spike_register[119] = spike119;        spike_register[120] = spike120;        spike_register[121] = spike121;        spike_register[122] = spike122;        spike_register[123] = spike123;        spike_register[124] = spike124;        spike_register[125] = spike125;        spike_register[126] = spike126;        spike_register[127] = spike127;        spike_register[128] = spike128;        spike_register[129] = spike129;        spike_register[130] = spike130;        spike_register[131] = spike131;        spike_register[132] = spike132;        spike_register[133] = spike133;        spike_register[134] = spike134;        spike_register[135] = spike135;        spike_register[136] = spike136;        spike_register[137] = spike137;        spike_register[138] = spike138;        spike_register[139] = spike139;        spike_register[140] = spike140;        spike_register[141] = spike141;        spike_register[142] = spike142;        spike_register[143] = spike143;        spike_register[144] = spike144;        spike_register[145] = spike145;        spike_register[146] = spike146;        spike_register[147] = spike147;        spike_register[148] = spike148;        spike_register[149] = spike149;
        #0.5
        if(clear == 1'b0) begin
            for(i3 = 100; i3 <=149; i3= i3+1) begin
                if(spike_register[i3] == 1 && lock3 == 0) begin
                    lock3 = 1;
                    for(j3 = connection_pointer[i3]; j3 < connection_pointer[i3+1]; j3= j3+1) begin
                        packet3 = #0.1 {neuron_addresses[i3], downstream_connections[j3]};
                    end
                    spike_register[i3] = 0;
                    lock3 = 0;
                end
            end
        end

    end
    always @(clear, lock4, spike150, spike151, spike152, spike153, spike154, spike155, spike156, spike157, spike158, spike159, spike160, spike161, spike162, spike163, spike164, spike165, spike166, spike167, spike168, spike169, spike170, spike171, spike172, spike173, spike174, spike175, spike176, spike177, spike178, spike179, spike180, spike181, spike182, spike183, spike184, spike185, spike186, spike187, spike188, spike189, spike190, spike191, spike192, spike193, spike194, spike195, spike196, spike197, spike198, spike199) begin
        spike_register[150] = spike150;        spike_register[151] = spike151;        spike_register[152] = spike152;        spike_register[153] = spike153;        spike_register[154] = spike154;        spike_register[155] = spike155;        spike_register[156] = spike156;        spike_register[157] = spike157;        spike_register[158] = spike158;        spike_register[159] = spike159;        spike_register[160] = spike160;        spike_register[161] = spike161;        spike_register[162] = spike162;        spike_register[163] = spike163;        spike_register[164] = spike164;        spike_register[165] = spike165;        spike_register[166] = spike166;        spike_register[167] = spike167;        spike_register[168] = spike168;        spike_register[169] = spike169;        spike_register[170] = spike170;        spike_register[171] = spike171;        spike_register[172] = spike172;        spike_register[173] = spike173;        spike_register[174] = spike174;        spike_register[175] = spike175;        spike_register[176] = spike176;        spike_register[177] = spike177;        spike_register[178] = spike178;        spike_register[179] = spike179;        spike_register[180] = spike180;        spike_register[181] = spike181;        spike_register[182] = spike182;        spike_register[183] = spike183;        spike_register[184] = spike184;        spike_register[185] = spike185;        spike_register[186] = spike186;        spike_register[187] = spike187;        spike_register[188] = spike188;        spike_register[189] = spike189;        spike_register[190] = spike190;        spike_register[191] = spike191;        spike_register[192] = spike192;        spike_register[193] = spike193;        spike_register[194] = spike194;        spike_register[195] = spike195;        spike_register[196] = spike196;        spike_register[197] = spike197;        spike_register[198] = spike198;        spike_register[199] = spike199;
        #0.5
        if(clear == 1'b0) begin
            for(i4 = 150; i4 <=199; i4= i4+1) begin
                if(spike_register[i4] == 1 && lock4 == 0) begin
                    lock4 = 1;
                    for(j4 = connection_pointer[i4]; j4 < connection_pointer[i4+1]; j4= j4+1) begin
                        packet4 = #0.1 {neuron_addresses[i4], downstream_connections[j4]};
                    end
                    spike_register[i4] = 0;
                    lock4 = 0;
                end
            end
        end

    end
    always @(clear, lock5, spike200, spike201, spike202, spike203, spike204, spike205, spike206, spike207, spike208, spike209, spike210, spike211, spike212, spike213, spike214, spike215, spike216, spike217, spike218, spike219, spike220, spike221, spike222, spike223, spike224, spike225, spike226, spike227, spike228, spike229, spike230, spike231, spike232, spike233, spike234, spike235, spike236, spike237, spike238, spike239, spike240, spike241, spike242, spike243, spike244, spike245, spike246, spike247, spike248, spike249) begin
        spike_register[200] = spike200;

        spike_register[201] = spike201;        spike_register[202] = spike202;        spike_register[203] = spike203;        spike_register[204] = spike204;        spike_register[205] = spike205;        spike_register[206] = spike206;        spike_register[207] = spike207;        spike_register[208] = spike208;        spike_register[209] = spike209;        spike_register[210] = spike210;        spike_register[211] = spike211;        spike_register[212] = spike212;        spike_register[213] = spike213;        spike_register[214] = spike214;        spike_register[215] = spike215;        spike_register[216] = spike216;        spike_register[217] = spike217;        spike_register[218] = spike218;        spike_register[219] = spike219;        spike_register[220] = spike220;        spike_register[221] = spike221;        spike_register[222] = spike222;        spike_register[223] = spike223;        spike_register[224] = spike224;        spike_register[225] = spike225;        spike_register[226] = spike226;        spike_register[227] = spike227;        spike_register[228] = spike228;        spike_register[229] = spike229;        spike_register[230] = spike230;        spike_register[231] = spike231;        spike_register[232] = spike232;        spike_register[233] = spike233;        spike_register[234] = spike234;        spike_register[235] = spike235;        spike_register[236] = spike236;        spike_register[237] = spike237;        spike_register[238] = spike238;        spike_register[239] = spike239;        spike_register[240] = spike240;        spike_register[241] = spike241;        spike_register[242] = spike242;        spike_register[243] = spike243;        spike_register[244] = spike244;        spike_register[245] = spike245;        spike_register[246] = spike246;        spike_register[247] = spike247;        spike_register[248] = spike248;        spike_register[249] = spike249;
        #0.5
        if(clear == 1'b0) begin
            for(i5 = 200; i5 <=249; i5= i5+1) begin
                if(spike_register[i5] == 1 && lock5 == 0) begin
                    lock5 = 1;
                    for(j5 = connection_pointer[i5]; j5 < connection_pointer[i5+1]; j5= j5+1) begin
                        packet5 = #0.1 {neuron_addresses[i5], downstream_connections[j5]};
                    end
                    spike_register[i5] = 0;
                    lock5 = 0;
                end
            end
        end

    end
    always @(clear, lock6, spike250, spike251, spike252, spike253, spike254, spike255, spike256, spike257, spike258, spike259, spike260, spike261, spike262, spike263, spike264, spike265, spike266, spike267, spike268, spike269, spike270, spike271, spike272, spike273, spike274, spike275, spike276, spike277, spike278, spike279, spike280, spike281, spike282, spike283, spike284, spike285, spike286, spike287, spike288, spike289, spike290, spike291, spike292, spike293, spike294, spike295, spike296, spike297, spike298, spike299) begin
        spike_register[250] = spike250;        spike_register[251] = spike251;        spike_register[252] = spike252;        spike_register[253] = spike253;        spike_register[254] = spike254;        spike_register[255] = spike255;        spike_register[256] = spike256;        spike_register[257] = spike257;        spike_register[258] = spike258;        spike_register[259] = spike259;        spike_register[260] = spike260;        spike_register[261] = spike261;        spike_register[262] = spike262;        spike_register[263] = spike263;        spike_register[264] = spike264;        spike_register[265] = spike265;        spike_register[266] = spike266;        spike_register[267] = spike267;        spike_register[268] = spike268;        spike_register[269] = spike269;        spike_register[270] = spike270;        spike_register[271] = spike271;        spike_register[272] = spike272;        spike_register[273] = spike273;        spike_register[274] = spike274;        spike_register[275] = spike275;        spike_register[276] = spike276;        spike_register[277] = spike277;        spike_register[278] = spike278;        spike_register[279] = spike279;        spike_register[280] = spike280;        spike_register[281] = spike281;        spike_register[282] = spike282;        spike_register[283] = spike283;        spike_register[284] = spike284;        spike_register[285] = spike285;        spike_register[286] = spike286;        spike_register[287] = spike287;        spike_register[288] = spike288;        spike_register[289] = spike289;        spike_register[290] = spike290;        spike_register[291] = spike291;        spike_register[292] = spike292;        spike_register[293] = spike293;        spike_register[294] = spike294;        spike_register[295] = spike295;        spike_register[296] = spike296;        spike_register[297] = spike297;        spike_register[298] = spike298;        spike_register[299] = spike299;
        #0.5
        if(clear == 1'b0) begin
            for(i6 = 250; i6 <=299; i6= i6+1) begin
                if(spike_register[i6] == 1 && lock6 == 0) begin
                    lock6 = 1;
                    for(j6 = connection_pointer[i6]; j6 < connection_pointer[i6+1]; j6= j6+1) begin
                        packet6 = #0.1 {neuron_addresses[i6], downstream_connections[j6]};
                    end
                    spike_register[i6] = 0;
                    lock6 = 0;
                end
            end
        end

    end
    always @(clear, lock7, spike300, spike301, spike302, spike303, spike304, spike305, spike306, spike307, spike308, spike309, spike310, spike311, spike312, spike313, spike314, spike315, spike316, spike317, spike318, spike319, spike320, spike321, spike322, spike323, spike324, spike325, spike326, spike327, spike328, spike329, spike330, spike331, spike332, spike333, spike334, spike335, spike336, spike337, spike338, spike339, spike340, spike341, spike342, spike343, spike344, spike345, spike346, spike347, spike348, spike349) begin
        spike_register[300] = spike300;

        spike_register[301] = spike301;        spike_register[302] = spike302;        spike_register[303] = spike303;        spike_register[304] = spike304;        spike_register[305] = spike305;        spike_register[306] = spike306;        spike_register[307] = spike307;        spike_register[308] = spike308;        spike_register[309] = spike309;        spike_register[310] = spike310;        spike_register[311] = spike311;        spike_register[312] = spike312;        spike_register[313] = spike313;        spike_register[314] = spike314;        spike_register[315] = spike315;        spike_register[316] = spike316;        spike_register[317] = spike317;        spike_register[318] = spike318;        spike_register[319] = spike319;        spike_register[320] = spike320;        spike_register[321] = spike321;        spike_register[322] = spike322;        spike_register[323] = spike323;        spike_register[324] = spike324;        spike_register[325] = spike325;        spike_register[326] = spike326;        spike_register[327] = spike327;        spike_register[328] = spike328;        spike_register[329] = spike329;        spike_register[330] = spike330;        spike_register[331] = spike331;        spike_register[332] = spike332;        spike_register[333] = spike333;        spike_register[334] = spike334;        spike_register[335] = spike335;        spike_register[336] = spike336;        spike_register[337] = spike337;        spike_register[338] = spike338;        spike_register[339] = spike339;        spike_register[340] = spike340;        spike_register[341] = spike341;        spike_register[342] = spike342;        spike_register[343] = spike343;        spike_register[344] = spike344;        spike_register[345] = spike345;        spike_register[346] = spike346;        spike_register[347] = spike347;        spike_register[348] = spike348;        spike_register[349] = spike349;
        #0.5
        if(clear == 1'b0) begin
            for(i7 = 300; i7 <=349; i7= i7+1) begin
                if(spike_register[i7] == 1 && lock7 == 0) begin
                    lock7 = 1;
                    for(j7 = connection_pointer[i7]; j7 < connection_pointer[i7+1]; j7= j7+1) begin
                        packet7 = #0.1 {neuron_addresses[i7], downstream_connections[j7]};
                    end
                    spike_register[i7] = 0;
                    lock7 = 0;
                end
            end
        end

    end
    always @(clear, lock8, spike350, spike351, spike352, spike353, spike354, spike355, spike356, spike357, spike358, spike359, spike360, spike361, spike362, spike363, spike364, spike365, spike366, spike367, spike368, spike369, spike370, spike371, spike372, spike373, spike374, spike375, spike376, spike377, spike378, spike379, spike380, spike381, spike382, spike383, spike384, spike385, spike386, spike387, spike388, spike389, spike390, spike391, spike392, spike393, spike394, spike395, spike396, spike397, spike398, spike399) begin
        spike_register[350] = spike350;        spike_register[351] = spike351;        spike_register[352] = spike352;        spike_register[353] = spike353;        spike_register[354] = spike354;        spike_register[355] = spike355;        spike_register[356] = spike356;        spike_register[357] = spike357;        spike_register[358] = spike358;        spike_register[359] = spike359;        spike_register[360] = spike360;        spike_register[361] = spike361;        spike_register[362] = spike362;        spike_register[363] = spike363;        spike_register[364] = spike364;        spike_register[365] = spike365;        spike_register[366] = spike366;        spike_register[367] = spike367;        spike_register[368] = spike368;        spike_register[369] = spike369;        spike_register[370] = spike370;        spike_register[371] = spike371;        spike_register[372] = spike372;        spike_register[373] = spike373;        spike_register[374] = spike374;        spike_register[375] = spike375;        spike_register[376] = spike376;        spike_register[377] = spike377;        spike_register[378] = spike378;        spike_register[379] = spike379;        spike_register[380] = spike380;        spike_register[381] = spike381;        spike_register[382] = spike382;        spike_register[383] = spike383;        spike_register[384] = spike384;        spike_register[385] = spike385;        spike_register[386] = spike386;        spike_register[387] = spike387;        spike_register[388] = spike388;        spike_register[389] = spike389;        spike_register[390] = spike390;        spike_register[391] = spike391;        spike_register[392] = spike392;        spike_register[393] = spike393;        spike_register[394] = spike394;        spike_register[395] = spike395;        spike_register[396] = spike396;        spike_register[397] = spike397;        spike_register[398] = spike398;        spike_register[399] = spike399;
        #0.5
        if(clear == 1'b0) begin
            for(i8 = 350; i8 <=399; i8= i8+1) begin
                if(spike_register[i8] == 1 && lock8 == 0) begin
                    lock8 = 1;
                    for(j8 = connection_pointer[i8]; j8 < connection_pointer[i8+1]; j8= j8+1) begin
                        packet8 = #0.1 {neuron_addresses[i8], downstream_connections[j8]};
                    end
                    spike_register[i8] = 0;
                    lock8 = 0;
                end
            end
        end

    end
    always @(clear, lock9, spike400, spike401, spike402, spike403, spike404, spike405, spike406, spike407, spike408, spike409, spike410, spike411, spike412, spike413, spike414, spike415, spike416, spike417, spike418, spike419, spike420, spike421, spike422, spike423, spike424, spike425, spike426, spike427, spike428, spike429, spike430, spike431, spike432, spike433, spike434, spike435, spike436, spike437, spike438, spike439, spike440, spike441, spike442, spike443, spike444, spike445, spike446, spike447, spike448, spike449) begin
        spike_register[400] = spike400;

        spike_register[401] = spike401;        spike_register[402] = spike402;        spike_register[403] = spike403;        spike_register[404] = spike404;        spike_register[405] = spike405;        spike_register[406] = spike406;        spike_register[407] = spike407;        spike_register[408] = spike408;        spike_register[409] = spike409;        spike_register[410] = spike410;        spike_register[411] = spike411;        spike_register[412] = spike412;        spike_register[413] = spike413;        spike_register[414] = spike414;        spike_register[415] = spike415;        spike_register[416] = spike416;        spike_register[417] = spike417;        spike_register[418] = spike418;        spike_register[419] = spike419;        spike_register[420] = spike420;        spike_register[421] = spike421;        spike_register[422] = spike422;        spike_register[423] = spike423;        spike_register[424] = spike424;        spike_register[425] = spike425;        spike_register[426] = spike426;        spike_register[427] = spike427;        spike_register[428] = spike428;        spike_register[429] = spike429;        spike_register[430] = spike430;        spike_register[431] = spike431;        spike_register[432] = spike432;        spike_register[433] = spike433;        spike_register[434] = spike434;        spike_register[435] = spike435;        spike_register[436] = spike436;        spike_register[437] = spike437;        spike_register[438] = spike438;        spike_register[439] = spike439;        spike_register[440] = spike440;        spike_register[441] = spike441;        spike_register[442] = spike442;        spike_register[443] = spike443;        spike_register[444] = spike444;        spike_register[445] = spike445;        spike_register[446] = spike446;        spike_register[447] = spike447;        spike_register[448] = spike448;        spike_register[449] = spike449;
        #0.5
        if(clear == 1'b0) begin
            for(i9 = 400; i9 <=449; i9= i9+1) begin
                if(spike_register[i9] == 1 && lock9 == 0) begin
                    lock9 = 1;
                    for(j9 = connection_pointer[i9]; j9 < connection_pointer[i9+1]; j9= j9+1) begin
                        packet9 = #0.1 {neuron_addresses[i9], downstream_connections[j9]};
                    end
                    spike_register[i9] = 0;
                    lock9 = 0;
                end
            end
        end

    end
    always @(clear, lock10, spike450, spike451, spike452, spike453, spike454, spike455, spike456, spike457, spike458, spike459, spike460, spike461, spike462, spike463, spike464, spike465, spike466, spike467, spike468, spike469, spike470, spike471, spike472, spike473, spike474, spike475, spike476, spike477, spike478, spike479, spike480, spike481, spike482, spike483, spike484, spike485, spike486, spike487, spike488, spike489, spike490, spike491, spike492, spike493, spike494, spike495, spike496, spike497, spike498, spike499) begin
        spike_register[450] = spike450;        spike_register[451] = spike451;        spike_register[452] = spike452;        spike_register[453] = spike453;        spike_register[454] = spike454;        spike_register[455] = spike455;        spike_register[456] = spike456;        spike_register[457] = spike457;        spike_register[458] = spike458;        spike_register[459] = spike459;        spike_register[460] = spike460;        spike_register[461] = spike461;        spike_register[462] = spike462;        spike_register[463] = spike463;        spike_register[464] = spike464;        spike_register[465] = spike465;        spike_register[466] = spike466;        spike_register[467] = spike467;        spike_register[468] = spike468;        spike_register[469] = spike469;        spike_register[470] = spike470;        spike_register[471] = spike471;        spike_register[472] = spike472;        spike_register[473] = spike473;        spike_register[474] = spike474;        spike_register[475] = spike475;        spike_register[476] = spike476;        spike_register[477] = spike477;        spike_register[478] = spike478;        spike_register[479] = spike479;        spike_register[480] = spike480;        spike_register[481] = spike481;        spike_register[482] = spike482;        spike_register[483] = spike483;        spike_register[484] = spike484;        spike_register[485] = spike485;        spike_register[486] = spike486;        spike_register[487] = spike487;        spike_register[488] = spike488;        spike_register[489] = spike489;        spike_register[490] = spike490;        spike_register[491] = spike491;        spike_register[492] = spike492;        spike_register[493] = spike493;        spike_register[494] = spike494;        spike_register[495] = spike495;        spike_register[496] = spike496;        spike_register[497] = spike497;        spike_register[498] = spike498;        spike_register[499] = spike499;
        #0.5
        if(clear == 1'b0) begin
            for(i10 = 450; i10 <=499; i10= i10+1) begin
                if(spike_register[i10] == 1 && lock10 == 0) begin
                    lock10 = 1;
                    for(j10 = connection_pointer[i10]; j10 < connection_pointer[i10+1]; j10= j10+1) begin
                        packet10 = #0.1 {neuron_addresses[i10], downstream_connections[j10]};
                    end
                    spike_register[i10] = 0;
                    lock10 = 0;
                end
            end
        end

    end
    always @(clear, lock11, spike500, spike501, spike502, spike503, spike504, spike505, spike506, spike507, spike508, spike509, spike510, spike511, spike512, spike513, spike514, spike515, spike516, spike517, spike518, spike519, spike520, spike521, spike522, spike523, spike524, spike525, spike526, spike527, spike528, spike529, spike530, spike531, spike532, spike533, spike534, spike535, spike536, spike537, spike538, spike539, spike540, spike541, spike542, spike543, spike544, spike545, spike546, spike547, spike548, spike549) begin
        spike_register[500] = spike500;

        spike_register[501] = spike501;        spike_register[502] = spike502;        spike_register[503] = spike503;        spike_register[504] = spike504;        spike_register[505] = spike505;        spike_register[506] = spike506;        spike_register[507] = spike507;        spike_register[508] = spike508;        spike_register[509] = spike509;        spike_register[510] = spike510;        spike_register[511] = spike511;        spike_register[512] = spike512;        spike_register[513] = spike513;        spike_register[514] = spike514;        spike_register[515] = spike515;        spike_register[516] = spike516;        spike_register[517] = spike517;        spike_register[518] = spike518;        spike_register[519] = spike519;        spike_register[520] = spike520;        spike_register[521] = spike521;        spike_register[522] = spike522;        spike_register[523] = spike523;        spike_register[524] = spike524;        spike_register[525] = spike525;        spike_register[526] = spike526;        spike_register[527] = spike527;        spike_register[528] = spike528;        spike_register[529] = spike529;        spike_register[530] = spike530;        spike_register[531] = spike531;        spike_register[532] = spike532;        spike_register[533] = spike533;        spike_register[534] = spike534;        spike_register[535] = spike535;        spike_register[536] = spike536;        spike_register[537] = spike537;        spike_register[538] = spike538;        spike_register[539] = spike539;        spike_register[540] = spike540;        spike_register[541] = spike541;        spike_register[542] = spike542;        spike_register[543] = spike543;        spike_register[544] = spike544;        spike_register[545] = spike545;        spike_register[546] = spike546;        spike_register[547] = spike547;        spike_register[548] = spike548;        spike_register[549] = spike549;
        #0.5
        if(clear == 1'b0) begin
            for(i11 = 500; i11 <=549; i11= i11+1) begin
                if(spike_register[i11] == 1 && lock11 == 0) begin
                    lock11 = 1;
                    for(j11 = connection_pointer[i11]; j11 < connection_pointer[i11+1]; j11= j11+1) begin
                        packet11 = #0.1 {neuron_addresses[i11], downstream_connections[j11]};
                    end
                    spike_register[i11] = 0;
                    lock11 = 0;
                end
            end
        end

    end
    always @(clear, lock12, spike550, spike551, spike552, spike553, spike554, spike555, spike556, spike557, spike558, spike559, spike560, spike561, spike562, spike563, spike564, spike565, spike566, spike567, spike568, spike569, spike570, spike571, spike572, spike573, spike574, spike575, spike576, spike577, spike578, spike579, spike580, spike581, spike582, spike583, spike584, spike585, spike586, spike587, spike588, spike589, spike590, spike591, spike592, spike593, spike594, spike595, spike596, spike597, spike598, spike599) begin
        spike_register[550] = spike550;        spike_register[551] = spike551;        spike_register[552] = spike552;        spike_register[553] = spike553;        spike_register[554] = spike554;        spike_register[555] = spike555;        spike_register[556] = spike556;        spike_register[557] = spike557;        spike_register[558] = spike558;        spike_register[559] = spike559;        spike_register[560] = spike560;        spike_register[561] = spike561;        spike_register[562] = spike562;        spike_register[563] = spike563;        spike_register[564] = spike564;        spike_register[565] = spike565;        spike_register[566] = spike566;        spike_register[567] = spike567;        spike_register[568] = spike568;        spike_register[569] = spike569;        spike_register[570] = spike570;        spike_register[571] = spike571;        spike_register[572] = spike572;        spike_register[573] = spike573;        spike_register[574] = spike574;        spike_register[575] = spike575;        spike_register[576] = spike576;        spike_register[577] = spike577;        spike_register[578] = spike578;        spike_register[579] = spike579;        spike_register[580] = spike580;        spike_register[581] = spike581;        spike_register[582] = spike582;        spike_register[583] = spike583;        spike_register[584] = spike584;        spike_register[585] = spike585;        spike_register[586] = spike586;        spike_register[587] = spike587;        spike_register[588] = spike588;        spike_register[589] = spike589;        spike_register[590] = spike590;        spike_register[591] = spike591;        spike_register[592] = spike592;        spike_register[593] = spike593;        spike_register[594] = spike594;        spike_register[595] = spike595;        spike_register[596] = spike596;        spike_register[597] = spike597;        spike_register[598] = spike598;        spike_register[599] = spike599;
        #0.5
        if(clear == 1'b0) begin
            for(i12 = 550; i12 <=599; i12= i12+1) begin
                if(spike_register[i12] == 1 && lock12 == 0) begin
                    lock12 = 1;
                    for(j12 = connection_pointer[i12]; j12 < connection_pointer[i12+1]; j12= j12+1) begin
                        packet12 = #0.1 {neuron_addresses[i12], downstream_connections[j12]};
                    end
                    spike_register[i12] = 0;
                    lock12 = 0;
                end
            end
        end

    end
    always @(clear, lock13, spike600, spike601, spike602, spike603, spike604, spike605, spike606, spike607, spike608, spike609, spike610, spike611, spike612, spike613, spike614, spike615, spike616, spike617, spike618, spike619, spike620, spike621, spike622, spike623, spike624, spike625, spike626, spike627, spike628, spike629, spike630, spike631, spike632, spike633, spike634, spike635, spike636, spike637, spike638, spike639, spike640, spike641, spike642, spike643, spike644, spike645, spike646, spike647, spike648, spike649) begin
        spike_register[600] = spike600;

        spike_register[601] = spike601;        spike_register[602] = spike602;        spike_register[603] = spike603;        spike_register[604] = spike604;        spike_register[605] = spike605;        spike_register[606] = spike606;        spike_register[607] = spike607;        spike_register[608] = spike608;        spike_register[609] = spike609;        spike_register[610] = spike610;        spike_register[611] = spike611;        spike_register[612] = spike612;        spike_register[613] = spike613;        spike_register[614] = spike614;        spike_register[615] = spike615;        spike_register[616] = spike616;        spike_register[617] = spike617;        spike_register[618] = spike618;        spike_register[619] = spike619;        spike_register[620] = spike620;        spike_register[621] = spike621;        spike_register[622] = spike622;        spike_register[623] = spike623;        spike_register[624] = spike624;        spike_register[625] = spike625;        spike_register[626] = spike626;        spike_register[627] = spike627;        spike_register[628] = spike628;        spike_register[629] = spike629;        spike_register[630] = spike630;        spike_register[631] = spike631;        spike_register[632] = spike632;        spike_register[633] = spike633;        spike_register[634] = spike634;        spike_register[635] = spike635;        spike_register[636] = spike636;        spike_register[637] = spike637;        spike_register[638] = spike638;        spike_register[639] = spike639;        spike_register[640] = spike640;        spike_register[641] = spike641;        spike_register[642] = spike642;        spike_register[643] = spike643;        spike_register[644] = spike644;        spike_register[645] = spike645;        spike_register[646] = spike646;        spike_register[647] = spike647;        spike_register[648] = spike648;        spike_register[649] = spike649;
        #0.5
        if(clear == 1'b0) begin
            for(i13 = 600; i13 <=649; i13= i13+1) begin
                if(spike_register[i13] == 1 && lock13 == 0) begin
                    lock13 = 1;
                    for(j13 = connection_pointer[i13]; j13 < connection_pointer[i13+1]; j13= j13+1) begin
                        packet13 = #0.1 {neuron_addresses[i13], downstream_connections[j13]};
                    end
                    spike_register[i13] = 0;
                    lock13 = 0;
                end
            end
        end

    end
    always @(clear, lock14, spike650, spike651, spike652, spike653, spike654, spike655, spike656, spike657, spike658, spike659, spike660, spike661, spike662, spike663, spike664, spike665, spike666, spike667, spike668, spike669, spike670, spike671, spike672, spike673, spike674, spike675, spike676, spike677, spike678, spike679, spike680, spike681, spike682, spike683, spike684, spike685, spike686, spike687, spike688, spike689, spike690, spike691, spike692, spike693, spike694, spike695, spike696, spike697, spike698, spike699) begin
        spike_register[650] = spike650;        spike_register[651] = spike651;        spike_register[652] = spike652;        spike_register[653] = spike653;        spike_register[654] = spike654;        spike_register[655] = spike655;        spike_register[656] = spike656;        spike_register[657] = spike657;        spike_register[658] = spike658;        spike_register[659] = spike659;        spike_register[660] = spike660;        spike_register[661] = spike661;        spike_register[662] = spike662;        spike_register[663] = spike663;        spike_register[664] = spike664;        spike_register[665] = spike665;        spike_register[666] = spike666;        spike_register[667] = spike667;        spike_register[668] = spike668;        spike_register[669] = spike669;        spike_register[670] = spike670;        spike_register[671] = spike671;        spike_register[672] = spike672;        spike_register[673] = spike673;        spike_register[674] = spike674;        spike_register[675] = spike675;        spike_register[676] = spike676;        spike_register[677] = spike677;        spike_register[678] = spike678;        spike_register[679] = spike679;        spike_register[680] = spike680;        spike_register[681] = spike681;        spike_register[682] = spike682;        spike_register[683] = spike683;        spike_register[684] = spike684;        spike_register[685] = spike685;        spike_register[686] = spike686;        spike_register[687] = spike687;        spike_register[688] = spike688;        spike_register[689] = spike689;        spike_register[690] = spike690;        spike_register[691] = spike691;        spike_register[692] = spike692;        spike_register[693] = spike693;        spike_register[694] = spike694;        spike_register[695] = spike695;        spike_register[696] = spike696;        spike_register[697] = spike697;        spike_register[698] = spike698;        spike_register[699] = spike699;
        #0.5
        if(clear == 1'b0) begin
            for(i14 = 650; i14 <=699; i14= i14+1) begin
                if(spike_register[i14] == 1 && lock14 == 0) begin
                    lock14 = 1;
                    for(j14 = connection_pointer[i14]; j14 < connection_pointer[i14+1]; j14= j14+1) begin
                        packet14 = #0.1 {neuron_addresses[i14], downstream_connections[j14]};
                    end
                    spike_register[i14] = 0;
                    lock14 = 0;
                end
            end
        end

    end
    always @(clear, lock15, spike700, spike701, spike702, spike703, spike704, spike705, spike706, spike707, spike708, spike709, spike710, spike711, spike712, spike713, spike714, spike715, spike716, spike717, spike718, spike719, spike720, spike721, spike722, spike723, spike724, spike725, spike726, spike727, spike728, spike729, spike730, spike731, spike732, spike733, spike734, spike735, spike736, spike737, spike738, spike739, spike740, spike741, spike742, spike743, spike744, spike745, spike746, spike747, spike748, spike749) begin
        spike_register[700] = spike700;

        spike_register[701] = spike701;        spike_register[702] = spike702;        spike_register[703] = spike703;        spike_register[704] = spike704;        spike_register[705] = spike705;        spike_register[706] = spike706;        spike_register[707] = spike707;        spike_register[708] = spike708;        spike_register[709] = spike709;        spike_register[710] = spike710;        spike_register[711] = spike711;        spike_register[712] = spike712;        spike_register[713] = spike713;        spike_register[714] = spike714;        spike_register[715] = spike715;        spike_register[716] = spike716;        spike_register[717] = spike717;        spike_register[718] = spike718;        spike_register[719] = spike719;        spike_register[720] = spike720;        spike_register[721] = spike721;        spike_register[722] = spike722;        spike_register[723] = spike723;        spike_register[724] = spike724;        spike_register[725] = spike725;        spike_register[726] = spike726;        spike_register[727] = spike727;        spike_register[728] = spike728;        spike_register[729] = spike729;        spike_register[730] = spike730;        spike_register[731] = spike731;        spike_register[732] = spike732;        spike_register[733] = spike733;        spike_register[734] = spike734;        spike_register[735] = spike735;        spike_register[736] = spike736;        spike_register[737] = spike737;        spike_register[738] = spike738;        spike_register[739] = spike739;        spike_register[740] = spike740;        spike_register[741] = spike741;        spike_register[742] = spike742;        spike_register[743] = spike743;        spike_register[744] = spike744;        spike_register[745] = spike745;        spike_register[746] = spike746;        spike_register[747] = spike747;        spike_register[748] = spike748;        spike_register[749] = spike749;
        #0.5
        if(clear == 1'b0) begin
            for(i15 = 700; i15 <=749; i15= i15+1) begin
                if(spike_register[i15] == 1 && lock15 == 0) begin
                    lock15 = 1;
                    for(j15 = connection_pointer[i15]; j15 < connection_pointer[i15+1]; j15= j15+1) begin
                        packet15 = #0.1 {neuron_addresses[i15], downstream_connections[j15]};
                    end
                    spike_register[i15] = 0;
                    lock15 = 0;
                end
            end
        end

    end
    always @(clear, lock16, spike750, spike751, spike752, spike753, spike754, spike755, spike756, spike757, spike758, spike759, spike760, spike761, spike762, spike763, spike764, spike765, spike766, spike767, spike768, spike769, spike770, spike771, spike772, spike773, spike774, spike775, spike776, spike777, spike778, spike779, spike780, spike781, spike782, spike783, spike784, spike785, spike786, spike787, spike788, spike789, spike790, spike791, spike792, spike793, spike794, spike795, spike796, spike797, spike798, spike799) begin
        spike_register[750] = spike750;        spike_register[751] = spike751;        spike_register[752] = spike752;        spike_register[753] = spike753;        spike_register[754] = spike754;        spike_register[755] = spike755;        spike_register[756] = spike756;        spike_register[757] = spike757;        spike_register[758] = spike758;        spike_register[759] = spike759;        spike_register[760] = spike760;        spike_register[761] = spike761;        spike_register[762] = spike762;        spike_register[763] = spike763;        spike_register[764] = spike764;        spike_register[765] = spike765;        spike_register[766] = spike766;        spike_register[767] = spike767;        spike_register[768] = spike768;        spike_register[769] = spike769;        spike_register[770] = spike770;        spike_register[771] = spike771;        spike_register[772] = spike772;        spike_register[773] = spike773;        spike_register[774] = spike774;        spike_register[775] = spike775;        spike_register[776] = spike776;        spike_register[777] = spike777;        spike_register[778] = spike778;        spike_register[779] = spike779;        spike_register[780] = spike780;        spike_register[781] = spike781;        spike_register[782] = spike782;        spike_register[783] = spike783;        spike_register[784] = spike784;        spike_register[785] = spike785;        spike_register[786] = spike786;        spike_register[787] = spike787;        spike_register[788] = spike788;        spike_register[789] = spike789;        spike_register[790] = spike790;        spike_register[791] = spike791;        spike_register[792] = spike792;        spike_register[793] = spike793;        spike_register[794] = spike794;        spike_register[795] = spike795;        spike_register[796] = spike796;        spike_register[797] = spike797;        spike_register[798] = spike798;        spike_register[799] = spike799;
        #0.5
        if(clear == 1'b0) begin
            for(i16 = 750; i16 <=799; i16= i16+1) begin
                if(spike_register[i16] == 1 && lock16 == 0) begin
                    lock16 = 1;
                    for(j16 = connection_pointer[i16]; j16 < connection_pointer[i16+1]; j16= j16+1) begin
                        packet16 = #0.1 {neuron_addresses[i16], downstream_connections[j16]};
                    end
                    spike_register[i16] = 0;
                    lock16 = 0;
                end
            end
        end

    end
    always @(clear, lock17, spike800, spike801, spike802, spike803, spike804, spike805, spike806, spike807, spike808, spike809, spike810, spike811, spike812, spike813, spike814, spike815, spike816, spike817, spike818, spike819, spike820, spike821, spike822, spike823, spike824, spike825, spike826, spike827, spike828, spike829, spike830, spike831, spike832, spike833, spike834, spike835, spike836, spike837, spike838, spike839, spike840, spike841, spike842, spike843, spike844, spike845, spike846, spike847, spike848, spike849) begin
        spike_register[800] = spike800;

        spike_register[801] = spike801;        spike_register[802] = spike802;        spike_register[803] = spike803;        spike_register[804] = spike804;        spike_register[805] = spike805;        spike_register[806] = spike806;        spike_register[807] = spike807;        spike_register[808] = spike808;        spike_register[809] = spike809;        spike_register[810] = spike810;        spike_register[811] = spike811;        spike_register[812] = spike812;        spike_register[813] = spike813;        spike_register[814] = spike814;        spike_register[815] = spike815;        spike_register[816] = spike816;        spike_register[817] = spike817;        spike_register[818] = spike818;        spike_register[819] = spike819;        spike_register[820] = spike820;        spike_register[821] = spike821;        spike_register[822] = spike822;        spike_register[823] = spike823;        spike_register[824] = spike824;        spike_register[825] = spike825;        spike_register[826] = spike826;        spike_register[827] = spike827;        spike_register[828] = spike828;        spike_register[829] = spike829;        spike_register[830] = spike830;        spike_register[831] = spike831;        spike_register[832] = spike832;        spike_register[833] = spike833;        spike_register[834] = spike834;        spike_register[835] = spike835;        spike_register[836] = spike836;        spike_register[837] = spike837;        spike_register[838] = spike838;        spike_register[839] = spike839;        spike_register[840] = spike840;        spike_register[841] = spike841;        spike_register[842] = spike842;        spike_register[843] = spike843;        spike_register[844] = spike844;        spike_register[845] = spike845;        spike_register[846] = spike846;        spike_register[847] = spike847;        spike_register[848] = spike848;        spike_register[849] = spike849;
        #0.5
        if(clear == 1'b0) begin
            for(i17 = 800; i17 <=849; i17= i17+1) begin
                if(spike_register[i17] == 1 && lock17 == 0) begin
                    lock17 = 1;
                    for(j17 = connection_pointer[i17]; j17 < connection_pointer[i17+1]; j17= j17+1) begin
                        packet17 = #0.1 {neuron_addresses[i17], downstream_connections[j17]};
                    end
                    spike_register[i17] = 0;
                    lock17 = 0;
                end
            end
        end

    end
    always @(clear, lock18, spike850, spike851, spike852, spike853, spike854, spike855, spike856, spike857, spike858, spike859, spike860, spike861, spike862, spike863, spike864, spike865, spike866, spike867, spike868, spike869, spike870, spike871, spike872, spike873, spike874, spike875, spike876, spike877, spike878, spike879, spike880, spike881, spike882, spike883, spike884, spike885, spike886, spike887, spike888, spike889, spike890, spike891, spike892, spike893, spike894, spike895, spike896, spike897, spike898, spike899) begin
        spike_register[850] = spike850;        spike_register[851] = spike851;        spike_register[852] = spike852;        spike_register[853] = spike853;        spike_register[854] = spike854;        spike_register[855] = spike855;        spike_register[856] = spike856;        spike_register[857] = spike857;        spike_register[858] = spike858;        spike_register[859] = spike859;        spike_register[860] = spike860;        spike_register[861] = spike861;        spike_register[862] = spike862;        spike_register[863] = spike863;        spike_register[864] = spike864;        spike_register[865] = spike865;        spike_register[866] = spike866;        spike_register[867] = spike867;        spike_register[868] = spike868;        spike_register[869] = spike869;        spike_register[870] = spike870;        spike_register[871] = spike871;        spike_register[872] = spike872;        spike_register[873] = spike873;        spike_register[874] = spike874;        spike_register[875] = spike875;        spike_register[876] = spike876;        spike_register[877] = spike877;        spike_register[878] = spike878;        spike_register[879] = spike879;        spike_register[880] = spike880;        spike_register[881] = spike881;        spike_register[882] = spike882;        spike_register[883] = spike883;        spike_register[884] = spike884;        spike_register[885] = spike885;        spike_register[886] = spike886;        spike_register[887] = spike887;        spike_register[888] = spike888;        spike_register[889] = spike889;        spike_register[890] = spike890;        spike_register[891] = spike891;        spike_register[892] = spike892;        spike_register[893] = spike893;        spike_register[894] = spike894;        spike_register[895] = spike895;        spike_register[896] = spike896;        spike_register[897] = spike897;        spike_register[898] = spike898;        spike_register[899] = spike899;
        #0.5
        if(clear == 1'b0) begin
            for(i18 = 850; i18 <=899; i18= i18+1) begin
                if(spike_register[i18] == 1 && lock18 == 0) begin
                    lock18 = 1;
                    for(j18 = connection_pointer[i18]; j18 < connection_pointer[i18+1]; j18= j18+1) begin
                        packet18 = #0.1 {neuron_addresses[i18], downstream_connections[j18]};
                    end
                    spike_register[i18] = 0;
                    lock18 = 0;
                end
            end
        end

    end
    always @(clear, lock19, spike900, spike901, spike902, spike903, spike904, spike905, spike906, spike907, spike908, spike909, spike910, spike911, spike912, spike913, spike914, spike915, spike916, spike917, spike918, spike919, spike920, spike921, spike922, spike923, spike924, spike925, spike926, spike927, spike928, spike929, spike930, spike931, spike932, spike933, spike934, spike935, spike936, spike937, spike938, spike939, spike940, spike941, spike942, spike943, spike944, spike945, spike946, spike947, spike948, spike949) begin
        spike_register[900] = spike900;

        spike_register[901] = spike901;        spike_register[902] = spike902;        spike_register[903] = spike903;        spike_register[904] = spike904;        spike_register[905] = spike905;        spike_register[906] = spike906;        spike_register[907] = spike907;        spike_register[908] = spike908;        spike_register[909] = spike909;        spike_register[910] = spike910;        spike_register[911] = spike911;        spike_register[912] = spike912;        spike_register[913] = spike913;        spike_register[914] = spike914;        spike_register[915] = spike915;        spike_register[916] = spike916;        spike_register[917] = spike917;        spike_register[918] = spike918;        spike_register[919] = spike919;        spike_register[920] = spike920;        spike_register[921] = spike921;        spike_register[922] = spike922;        spike_register[923] = spike923;        spike_register[924] = spike924;        spike_register[925] = spike925;        spike_register[926] = spike926;        spike_register[927] = spike927;        spike_register[928] = spike928;        spike_register[929] = spike929;        spike_register[930] = spike930;        spike_register[931] = spike931;        spike_register[932] = spike932;        spike_register[933] = spike933;        spike_register[934] = spike934;        spike_register[935] = spike935;        spike_register[936] = spike936;        spike_register[937] = spike937;        spike_register[938] = spike938;        spike_register[939] = spike939;        spike_register[940] = spike940;        spike_register[941] = spike941;        spike_register[942] = spike942;        spike_register[943] = spike943;        spike_register[944] = spike944;        spike_register[945] = spike945;        spike_register[946] = spike946;        spike_register[947] = spike947;        spike_register[948] = spike948;        spike_register[949] = spike949;
        #0.5
        if(clear == 1'b0) begin
            for(i19 = 900; i19 <=949; i19= i19+1) begin
                if(spike_register[i19] == 1 && lock19 == 0) begin
                    lock19 = 1;
                    for(j19 = connection_pointer[i19]; j19 < connection_pointer[i19+1]; j19= j19+1) begin
                        packet19 = #0.1 {neuron_addresses[i19], downstream_connections[j19]};
                    end
                    spike_register[i19] = 0;
                    lock19 = 0;
                end
            end
        end

    end
    always @(clear, lock20, spike950, spike951, spike952, spike953, spike954, spike955, spike956, spike957, spike958, spike959, spike960, spike961, spike962, spike963, spike964, spike965, spike966, spike967, spike968, spike969, spike970, spike971, spike972, spike973, spike974, spike975, spike976, spike977, spike978, spike979, spike980, spike981, spike982, spike983, spike984, spike985, spike986, spike987, spike988, spike989, spike990, spike991, spike992, spike993, spike994, spike995, spike996, spike997, spike998, spike999) begin
        spike_register[950] = spike950;        spike_register[951] = spike951;        spike_register[952] = spike952;        spike_register[953] = spike953;        spike_register[954] = spike954;        spike_register[955] = spike955;        spike_register[956] = spike956;        spike_register[957] = spike957;        spike_register[958] = spike958;        spike_register[959] = spike959;        spike_register[960] = spike960;        spike_register[961] = spike961;        spike_register[962] = spike962;        spike_register[963] = spike963;        spike_register[964] = spike964;        spike_register[965] = spike965;        spike_register[966] = spike966;        spike_register[967] = spike967;        spike_register[968] = spike968;        spike_register[969] = spike969;        spike_register[970] = spike970;        spike_register[971] = spike971;        spike_register[972] = spike972;        spike_register[973] = spike973;        spike_register[974] = spike974;        spike_register[975] = spike975;        spike_register[976] = spike976;        spike_register[977] = spike977;        spike_register[978] = spike978;        spike_register[979] = spike979;        spike_register[980] = spike980;        spike_register[981] = spike981;        spike_register[982] = spike982;        spike_register[983] = spike983;        spike_register[984] = spike984;        spike_register[985] = spike985;        spike_register[986] = spike986;        spike_register[987] = spike987;        spike_register[988] = spike988;        spike_register[989] = spike989;        spike_register[990] = spike990;        spike_register[991] = spike991;        spike_register[992] = spike992;        spike_register[993] = spike993;        spike_register[994] = spike994;        spike_register[995] = spike995;        spike_register[996] = spike996;        spike_register[997] = spike997;        spike_register[998] = spike998;        spike_register[999] = spike999;
        #0.5
        if(clear == 1'b0) begin
            for(i20 = 950; i20 <=999; i20= i20+1) begin
                if(spike_register[i20] == 1 && lock20 == 0) begin
                    lock20 = 1;
                    for(j20 = connection_pointer[i20]; j20 < connection_pointer[i20+1]; j20= j20+1) begin
                        packet20 = #0.1 {neuron_addresses[i20], downstream_connections[j20]};
                    end
                    spike_register[i20] = 0;
                    lock20 = 0;
                end
            end
        end

    end
    always @(clear, lock21, spike1000, spike1001, spike1002, spike1003, spike1004, spike1005, spike1006, spike1007, spike1008, spike1009, spike1010, spike1011, spike1012, spike1013, spike1014, spike1015, spike1016, spike1017, spike1018, spike1019, spike1020, spike1021, spike1022, spike1023) begin
        spike_register[1000] = spike1000;

        spike_register[1001] = spike1001;        spike_register[1002] = spike1002;        spike_register[1003] = spike1003;        spike_register[1004] = spike1004;        spike_register[1005] = spike1005;        spike_register[1006] = spike1006;        spike_register[1007] = spike1007;        spike_register[1008] = spike1008;        spike_register[1009] = spike1009;        spike_register[1010] = spike1010;        spike_register[1011] = spike1011;        spike_register[1012] = spike1012;        spike_register[1013] = spike1013;        spike_register[1014] = spike1014;        spike_register[1015] = spike1015;        spike_register[1016] = spike1016;        spike_register[1017] = spike1017;        spike_register[1018] = spike1018;        spike_register[1019] = spike1019;        spike_register[1020] = spike1020;        spike_register[1021] = spike1021;        spike_register[1022] = spike1022;        spike_register[1023] = spike1023;
        #0.5
        if(clear == 1'b0) begin
            for(i21 = 1000; i21 <=1049; i21= i21+1) begin
                if(spike_register[i21] == 1 && lock21 == 0) begin
                    lock21 = 1;
                    for(j21 = connection_pointer[i21]; j21 < connection_pointer[i21+1]; j21= j21+1) begin
                        packet21 = #0.1 {neuron_addresses[i21], downstream_connections[j21]};
                    end
                    spike_register[i21] = 0;
                    lock21 = 0;
                end
            end
        end

    end
    always @(packet1) begin 
        spike_origin = packet1[23:12];
        spike_destination = packet1[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet2) begin 
        spike_origin = packet2[23:12];
        spike_destination = packet2[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet3) begin 
        spike_origin = packet3[23:12];
        spike_destination = packet3[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet4) begin 
        spike_origin = packet4[23:12];
        spike_destination = packet4[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet5) begin 
        spike_origin = packet5[23:12];
        spike_destination = packet5[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet6) begin 
        spike_origin = packet6[23:12];
        spike_destination = packet6[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet7) begin 
        spike_origin = packet7[23:12];
        spike_destination = packet7[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet8) begin 
        spike_origin = packet8[23:12];
        spike_destination = packet8[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet9) begin 
        spike_origin = packet9[23:12];
        spike_destination = packet9[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet10) begin 
        spike_origin = packet10[23:12];
        spike_destination = packet10[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet11) begin 
        spike_origin = packet11[23:12];
        spike_destination = packet11[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet12) begin 
        spike_origin = packet12[23:12];
        spike_destination = packet12[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet13) begin 
        spike_origin = packet13[23:12];
        spike_destination = packet13[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet14) begin 
        spike_origin = packet14[23:12];
        spike_destination = packet14[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet15) begin 
        spike_origin = packet15[23:12];
        spike_destination = packet15[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet16) begin 
        spike_origin = packet16[23:12];
        spike_destination = packet16[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet17) begin 
        spike_origin = packet17[23:12];
        spike_destination = packet17[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet18) begin 
        spike_origin = packet18[23:12];
        spike_destination = packet18[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet19) begin 
        spike_origin = packet19[23:12];
        spike_destination = packet19[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet20) begin 
        spike_origin = packet20[23:12];
        spike_destination = packet20[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet21) begin 
        spike_origin = packet21[23:12];
        spike_destination = packet21[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(spike_out_source_array[0]) begin 
        spike_out_source0 = spike_out_source_array[0];
    end
    always @(spike_out_source_array[1]) begin 
        spike_out_source1 = spike_out_source_array[1];
    end
    always @(spike_out_source_array[2]) begin 
        spike_out_source2 = spike_out_source_array[2];
    end
    always @(spike_out_source_array[3]) begin 
        spike_out_source3 = spike_out_source_array[3];
    end
    always @(spike_out_source_array[4]) begin 
        spike_out_source4 = spike_out_source_array[4];
    end
    always @(spike_out_source_array[5]) begin 
        spike_out_source5 = spike_out_source_array[5];
    end
    always @(spike_out_source_array[6]) begin 
        spike_out_source6 = spike_out_source_array[6];
    end
    always @(spike_out_source_array[7]) begin 
        spike_out_source7 = spike_out_source_array[7];
    end
    always @(spike_out_source_array[8]) begin 
        spike_out_source8 = spike_out_source_array[8];
    end
    always @(spike_out_source_array[9]) begin 
        spike_out_source9 = spike_out_source_array[9];
    end
    always @(spike_out_source_array[10]) begin 
        spike_out_source10 = spike_out_source_array[10];
    end
    always @(spike_out_source_array[11]) begin 
        spike_out_source11 = spike_out_source_array[11];
    end
    always @(spike_out_source_array[12]) begin 
        spike_out_source12 = spike_out_source_array[12];
    end
    always @(spike_out_source_array[13]) begin 
        spike_out_source13 = spike_out_source_array[13];
    end
    always @(spike_out_source_array[14]) begin 
        spike_out_source14 = spike_out_source_array[14];
    end
    always @(spike_out_source_array[15]) begin 
        spike_out_source15 = spike_out_source_array[15];
    end
    always @(spike_out_source_array[16]) begin 
        spike_out_source16 = spike_out_source_array[16];
    end
    always @(spike_out_source_array[17]) begin 
        spike_out_source17 = spike_out_source_array[17];
    end
    always @(spike_out_source_array[18]) begin 
        spike_out_source18 = spike_out_source_array[18];
    end
    always @(spike_out_source_array[19]) begin 
        spike_out_source19 = spike_out_source_array[19];
    end
    always @(spike_out_source_array[20]) begin 
        spike_out_source20 = spike_out_source_array[20];
    end
    always @(spike_out_source_array[21]) begin 
        spike_out_source21 = spike_out_source_array[21];
    end
    always @(spike_out_source_array[22]) begin 
        spike_out_source22 = spike_out_source_array[22];
    end
    always @(spike_out_source_array[23]) begin 
        spike_out_source23 = spike_out_source_array[23];
    end
    always @(spike_out_source_array[24]) begin 
        spike_out_source24 = spike_out_source_array[24];
    end
    always @(spike_out_source_array[25]) begin 
        spike_out_source25 = spike_out_source_array[25];
    end
    always @(spike_out_source_array[26]) begin 
        spike_out_source26 = spike_out_source_array[26];
    end
    always @(spike_out_source_array[27]) begin 
        spike_out_source27 = spike_out_source_array[27];
    end
    always @(spike_out_source_array[28]) begin 
        spike_out_source28 = spike_out_source_array[28];
    end
    always @(spike_out_source_array[29]) begin 
        spike_out_source29 = spike_out_source_array[29];
    end
    always @(spike_out_source_array[30]) begin 
        spike_out_source30 = spike_out_source_array[30];
    end
    always @(spike_out_source_array[31]) begin 
        spike_out_source31 = spike_out_source_array[31];
    end
    always @(spike_out_source_array[32]) begin 
        spike_out_source32 = spike_out_source_array[32];
    end
    always @(spike_out_source_array[33]) begin 
        spike_out_source33 = spike_out_source_array[33];
    end
    always @(spike_out_source_array[34]) begin 
        spike_out_source34 = spike_out_source_array[34];
    end
    always @(spike_out_source_array[35]) begin 
        spike_out_source35 = spike_out_source_array[35];
    end
    always @(spike_out_source_array[36]) begin 
        spike_out_source36 = spike_out_source_array[36];
    end
    always @(spike_out_source_array[37]) begin 
        spike_out_source37 = spike_out_source_array[37];
    end
    always @(spike_out_source_array[38]) begin 
        spike_out_source38 = spike_out_source_array[38];
    end
    always @(spike_out_source_array[39]) begin 
        spike_out_source39 = spike_out_source_array[39];
    end
    always @(spike_out_source_array[40]) begin 
        spike_out_source40 = spike_out_source_array[40];
    end
    always @(spike_out_source_array[41]) begin 
        spike_out_source41 = spike_out_source_array[41];
    end
    always @(spike_out_source_array[42]) begin 
        spike_out_source42 = spike_out_source_array[42];
    end
    always @(spike_out_source_array[43]) begin 
        spike_out_source43 = spike_out_source_array[43];
    end
    always @(spike_out_source_array[44]) begin 
        spike_out_source44 = spike_out_source_array[44];
    end
    always @(spike_out_source_array[45]) begin 
        spike_out_source45 = spike_out_source_array[45];
    end
    always @(spike_out_source_array[46]) begin 
        spike_out_source46 = spike_out_source_array[46];
    end
    always @(spike_out_source_array[47]) begin 
        spike_out_source47 = spike_out_source_array[47];
    end
    always @(spike_out_source_array[48]) begin 
        spike_out_source48 = spike_out_source_array[48];
    end
    always @(spike_out_source_array[49]) begin 
        spike_out_source49 = spike_out_source_array[49];
    end
    always @(spike_out_source_array[50]) begin 
        spike_out_source50 = spike_out_source_array[50];
    end
    always @(spike_out_source_array[51]) begin 
        spike_out_source51 = spike_out_source_array[51];
    end
    always @(spike_out_source_array[52]) begin 
        spike_out_source52 = spike_out_source_array[52];
    end
    always @(spike_out_source_array[53]) begin 
        spike_out_source53 = spike_out_source_array[53];
    end
    always @(spike_out_source_array[54]) begin 
        spike_out_source54 = spike_out_source_array[54];
    end
    always @(spike_out_source_array[55]) begin 
        spike_out_source55 = spike_out_source_array[55];
    end
    always @(spike_out_source_array[56]) begin 
        spike_out_source56 = spike_out_source_array[56];
    end
    always @(spike_out_source_array[57]) begin 
        spike_out_source57 = spike_out_source_array[57];
    end
    always @(spike_out_source_array[58]) begin 
        spike_out_source58 = spike_out_source_array[58];
    end
    always @(spike_out_source_array[59]) begin 
        spike_out_source59 = spike_out_source_array[59];
    end
    always @(spike_out_source_array[60]) begin 
        spike_out_source60 = spike_out_source_array[60];
    end
    always @(spike_out_source_array[61]) begin 
        spike_out_source61 = spike_out_source_array[61];
    end
    always @(spike_out_source_array[62]) begin 
        spike_out_source62 = spike_out_source_array[62];
    end
    always @(spike_out_source_array[63]) begin 
        spike_out_source63 = spike_out_source_array[63];
    end
    always @(spike_out_source_array[64]) begin 
        spike_out_source64 = spike_out_source_array[64];
    end
    always @(spike_out_source_array[65]) begin 
        spike_out_source65 = spike_out_source_array[65];
    end
    always @(spike_out_source_array[66]) begin 
        spike_out_source66 = spike_out_source_array[66];
    end
    always @(spike_out_source_array[67]) begin 
        spike_out_source67 = spike_out_source_array[67];
    end
    always @(spike_out_source_array[68]) begin 
        spike_out_source68 = spike_out_source_array[68];
    end
    always @(spike_out_source_array[69]) begin 
        spike_out_source69 = spike_out_source_array[69];
    end
    always @(spike_out_source_array[70]) begin 
        spike_out_source70 = spike_out_source_array[70];
    end
    always @(spike_out_source_array[71]) begin 
        spike_out_source71 = spike_out_source_array[71];
    end
    always @(spike_out_source_array[72]) begin 
        spike_out_source72 = spike_out_source_array[72];
    end
    always @(spike_out_source_array[73]) begin 
        spike_out_source73 = spike_out_source_array[73];
    end
    always @(spike_out_source_array[74]) begin 
        spike_out_source74 = spike_out_source_array[74];
    end
    always @(spike_out_source_array[75]) begin 
        spike_out_source75 = spike_out_source_array[75];
    end
    always @(spike_out_source_array[76]) begin 
        spike_out_source76 = spike_out_source_array[76];
    end
    always @(spike_out_source_array[77]) begin 
        spike_out_source77 = spike_out_source_array[77];
    end
    always @(spike_out_source_array[78]) begin 
        spike_out_source78 = spike_out_source_array[78];
    end
    always @(spike_out_source_array[79]) begin 
        spike_out_source79 = spike_out_source_array[79];
    end
    always @(spike_out_source_array[80]) begin 
        spike_out_source80 = spike_out_source_array[80];
    end
    always @(spike_out_source_array[81]) begin 
        spike_out_source81 = spike_out_source_array[81];
    end
    always @(spike_out_source_array[82]) begin 
        spike_out_source82 = spike_out_source_array[82];
    end
    always @(spike_out_source_array[83]) begin 
        spike_out_source83 = spike_out_source_array[83];
    end
    always @(spike_out_source_array[84]) begin 
        spike_out_source84 = spike_out_source_array[84];
    end
    always @(spike_out_source_array[85]) begin 
        spike_out_source85 = spike_out_source_array[85];
    end
    always @(spike_out_source_array[86]) begin 
        spike_out_source86 = spike_out_source_array[86];
    end
    always @(spike_out_source_array[87]) begin 
        spike_out_source87 = spike_out_source_array[87];
    end
    always @(spike_out_source_array[88]) begin 
        spike_out_source88 = spike_out_source_array[88];
    end
    always @(spike_out_source_array[89]) begin 
        spike_out_source89 = spike_out_source_array[89];
    end
    always @(spike_out_source_array[90]) begin 
        spike_out_source90 = spike_out_source_array[90];
    end
    always @(spike_out_source_array[91]) begin 
        spike_out_source91 = spike_out_source_array[91];
    end
    always @(spike_out_source_array[92]) begin 
        spike_out_source92 = spike_out_source_array[92];
    end
    always @(spike_out_source_array[93]) begin 
        spike_out_source93 = spike_out_source_array[93];
    end
    always @(spike_out_source_array[94]) begin 
        spike_out_source94 = spike_out_source_array[94];
    end
    always @(spike_out_source_array[95]) begin 
        spike_out_source95 = spike_out_source_array[95];
    end
    always @(spike_out_source_array[96]) begin 
        spike_out_source96 = spike_out_source_array[96];
    end
    always @(spike_out_source_array[97]) begin 
        spike_out_source97 = spike_out_source_array[97];
    end
    always @(spike_out_source_array[98]) begin 
        spike_out_source98 = spike_out_source_array[98];
    end
    always @(spike_out_source_array[99]) begin 
        spike_out_source99 = spike_out_source_array[99];
    end
    always @(spike_out_source_array[100]) begin 
        spike_out_source100 = spike_out_source_array[100];
    end
    always @(spike_out_source_array[101]) begin 
        spike_out_source101 = spike_out_source_array[101];
    end
    always @(spike_out_source_array[102]) begin 
        spike_out_source102 = spike_out_source_array[102];
    end
    always @(spike_out_source_array[103]) begin 
        spike_out_source103 = spike_out_source_array[103];
    end
    always @(spike_out_source_array[104]) begin 
        spike_out_source104 = spike_out_source_array[104];
    end
    always @(spike_out_source_array[105]) begin 
        spike_out_source105 = spike_out_source_array[105];
    end
    always @(spike_out_source_array[106]) begin 
        spike_out_source106 = spike_out_source_array[106];
    end
    always @(spike_out_source_array[107]) begin 
        spike_out_source107 = spike_out_source_array[107];
    end
    always @(spike_out_source_array[108]) begin 
        spike_out_source108 = spike_out_source_array[108];
    end
    always @(spike_out_source_array[109]) begin 
        spike_out_source109 = spike_out_source_array[109];
    end
    always @(spike_out_source_array[110]) begin 
        spike_out_source110 = spike_out_source_array[110];
    end
    always @(spike_out_source_array[111]) begin 
        spike_out_source111 = spike_out_source_array[111];
    end
    always @(spike_out_source_array[112]) begin 
        spike_out_source112 = spike_out_source_array[112];
    end
    always @(spike_out_source_array[113]) begin 
        spike_out_source113 = spike_out_source_array[113];
    end
    always @(spike_out_source_array[114]) begin 
        spike_out_source114 = spike_out_source_array[114];
    end
    always @(spike_out_source_array[115]) begin 
        spike_out_source115 = spike_out_source_array[115];
    end
    always @(spike_out_source_array[116]) begin 
        spike_out_source116 = spike_out_source_array[116];
    end
    always @(spike_out_source_array[117]) begin 
        spike_out_source117 = spike_out_source_array[117];
    end
    always @(spike_out_source_array[118]) begin 
        spike_out_source118 = spike_out_source_array[118];
    end
    always @(spike_out_source_array[119]) begin 
        spike_out_source119 = spike_out_source_array[119];
    end
    always @(spike_out_source_array[120]) begin 
        spike_out_source120 = spike_out_source_array[120];
    end
    always @(spike_out_source_array[121]) begin 
        spike_out_source121 = spike_out_source_array[121];
    end
    always @(spike_out_source_array[122]) begin 
        spike_out_source122 = spike_out_source_array[122];
    end
    always @(spike_out_source_array[123]) begin 
        spike_out_source123 = spike_out_source_array[123];
    end
    always @(spike_out_source_array[124]) begin 
        spike_out_source124 = spike_out_source_array[124];
    end
    always @(spike_out_source_array[125]) begin 
        spike_out_source125 = spike_out_source_array[125];
    end
    always @(spike_out_source_array[126]) begin 
        spike_out_source126 = spike_out_source_array[126];
    end
    always @(spike_out_source_array[127]) begin 
        spike_out_source127 = spike_out_source_array[127];
    end
    always @(spike_out_source_array[128]) begin 
        spike_out_source128 = spike_out_source_array[128];
    end
    always @(spike_out_source_array[129]) begin 
        spike_out_source129 = spike_out_source_array[129];
    end
    always @(spike_out_source_array[130]) begin 
        spike_out_source130 = spike_out_source_array[130];
    end
    always @(spike_out_source_array[131]) begin 
        spike_out_source131 = spike_out_source_array[131];
    end
    always @(spike_out_source_array[132]) begin 
        spike_out_source132 = spike_out_source_array[132];
    end
    always @(spike_out_source_array[133]) begin 
        spike_out_source133 = spike_out_source_array[133];
    end
    always @(spike_out_source_array[134]) begin 
        spike_out_source134 = spike_out_source_array[134];
    end
    always @(spike_out_source_array[135]) begin 
        spike_out_source135 = spike_out_source_array[135];
    end
    always @(spike_out_source_array[136]) begin 
        spike_out_source136 = spike_out_source_array[136];
    end
    always @(spike_out_source_array[137]) begin 
        spike_out_source137 = spike_out_source_array[137];
    end
    always @(spike_out_source_array[138]) begin 
        spike_out_source138 = spike_out_source_array[138];
    end
    always @(spike_out_source_array[139]) begin 
        spike_out_source139 = spike_out_source_array[139];
    end
    always @(spike_out_source_array[140]) begin 
        spike_out_source140 = spike_out_source_array[140];
    end
    always @(spike_out_source_array[141]) begin 
        spike_out_source141 = spike_out_source_array[141];
    end
    always @(spike_out_source_array[142]) begin 
        spike_out_source142 = spike_out_source_array[142];
    end
    always @(spike_out_source_array[143]) begin 
        spike_out_source143 = spike_out_source_array[143];
    end
    always @(spike_out_source_array[144]) begin 
        spike_out_source144 = spike_out_source_array[144];
    end
    always @(spike_out_source_array[145]) begin 
        spike_out_source145 = spike_out_source_array[145];
    end
    always @(spike_out_source_array[146]) begin 
        spike_out_source146 = spike_out_source_array[146];
    end
    always @(spike_out_source_array[147]) begin 
        spike_out_source147 = spike_out_source_array[147];
    end
    always @(spike_out_source_array[148]) begin 
        spike_out_source148 = spike_out_source_array[148];
    end
    always @(spike_out_source_array[149]) begin 
        spike_out_source149 = spike_out_source_array[149];
    end
    always @(spike_out_source_array[150]) begin 
        spike_out_source150 = spike_out_source_array[150];
    end
    always @(spike_out_source_array[151]) begin 
        spike_out_source151 = spike_out_source_array[151];
    end
    always @(spike_out_source_array[152]) begin 
        spike_out_source152 = spike_out_source_array[152];
    end
    always @(spike_out_source_array[153]) begin 
        spike_out_source153 = spike_out_source_array[153];
    end
    always @(spike_out_source_array[154]) begin 
        spike_out_source154 = spike_out_source_array[154];
    end
    always @(spike_out_source_array[155]) begin 
        spike_out_source155 = spike_out_source_array[155];
    end
    always @(spike_out_source_array[156]) begin 
        spike_out_source156 = spike_out_source_array[156];
    end
    always @(spike_out_source_array[157]) begin 
        spike_out_source157 = spike_out_source_array[157];
    end
    always @(spike_out_source_array[158]) begin 
        spike_out_source158 = spike_out_source_array[158];
    end
    always @(spike_out_source_array[159]) begin 
        spike_out_source159 = spike_out_source_array[159];
    end
    always @(spike_out_source_array[160]) begin 
        spike_out_source160 = spike_out_source_array[160];
    end
    always @(spike_out_source_array[161]) begin 
        spike_out_source161 = spike_out_source_array[161];
    end
    always @(spike_out_source_array[162]) begin 
        spike_out_source162 = spike_out_source_array[162];
    end
    always @(spike_out_source_array[163]) begin 
        spike_out_source163 = spike_out_source_array[163];
    end
    always @(spike_out_source_array[164]) begin 
        spike_out_source164 = spike_out_source_array[164];
    end
    always @(spike_out_source_array[165]) begin 
        spike_out_source165 = spike_out_source_array[165];
    end
    always @(spike_out_source_array[166]) begin 
        spike_out_source166 = spike_out_source_array[166];
    end
    always @(spike_out_source_array[167]) begin 
        spike_out_source167 = spike_out_source_array[167];
    end
    always @(spike_out_source_array[168]) begin 
        spike_out_source168 = spike_out_source_array[168];
    end
    always @(spike_out_source_array[169]) begin 
        spike_out_source169 = spike_out_source_array[169];
    end
    always @(spike_out_source_array[170]) begin 
        spike_out_source170 = spike_out_source_array[170];
    end
    always @(spike_out_source_array[171]) begin 
        spike_out_source171 = spike_out_source_array[171];
    end
    always @(spike_out_source_array[172]) begin 
        spike_out_source172 = spike_out_source_array[172];
    end
    always @(spike_out_source_array[173]) begin 
        spike_out_source173 = spike_out_source_array[173];
    end
    always @(spike_out_source_array[174]) begin 
        spike_out_source174 = spike_out_source_array[174];
    end
    always @(spike_out_source_array[175]) begin 
        spike_out_source175 = spike_out_source_array[175];
    end
    always @(spike_out_source_array[176]) begin 
        spike_out_source176 = spike_out_source_array[176];
    end
    always @(spike_out_source_array[177]) begin 
        spike_out_source177 = spike_out_source_array[177];
    end
    always @(spike_out_source_array[178]) begin 
        spike_out_source178 = spike_out_source_array[178];
    end
    always @(spike_out_source_array[179]) begin 
        spike_out_source179 = spike_out_source_array[179];
    end
    always @(spike_out_source_array[180]) begin 
        spike_out_source180 = spike_out_source_array[180];
    end
    always @(spike_out_source_array[181]) begin 
        spike_out_source181 = spike_out_source_array[181];
    end
    always @(spike_out_source_array[182]) begin 
        spike_out_source182 = spike_out_source_array[182];
    end
    always @(spike_out_source_array[183]) begin 
        spike_out_source183 = spike_out_source_array[183];
    end
    always @(spike_out_source_array[184]) begin 
        spike_out_source184 = spike_out_source_array[184];
    end
    always @(spike_out_source_array[185]) begin 
        spike_out_source185 = spike_out_source_array[185];
    end
    always @(spike_out_source_array[186]) begin 
        spike_out_source186 = spike_out_source_array[186];
    end
    always @(spike_out_source_array[187]) begin 
        spike_out_source187 = spike_out_source_array[187];
    end
    always @(spike_out_source_array[188]) begin 
        spike_out_source188 = spike_out_source_array[188];
    end
    always @(spike_out_source_array[189]) begin 
        spike_out_source189 = spike_out_source_array[189];
    end
    always @(spike_out_source_array[190]) begin 
        spike_out_source190 = spike_out_source_array[190];
    end
    always @(spike_out_source_array[191]) begin 
        spike_out_source191 = spike_out_source_array[191];
    end
    always @(spike_out_source_array[192]) begin 
        spike_out_source192 = spike_out_source_array[192];
    end
    always @(spike_out_source_array[193]) begin 
        spike_out_source193 = spike_out_source_array[193];
    end
    always @(spike_out_source_array[194]) begin 
        spike_out_source194 = spike_out_source_array[194];
    end
    always @(spike_out_source_array[195]) begin 
        spike_out_source195 = spike_out_source_array[195];
    end
    always @(spike_out_source_array[196]) begin 
        spike_out_source196 = spike_out_source_array[196];
    end
    always @(spike_out_source_array[197]) begin 
        spike_out_source197 = spike_out_source_array[197];
    end
    always @(spike_out_source_array[198]) begin 
        spike_out_source198 = spike_out_source_array[198];
    end
    always @(spike_out_source_array[199]) begin 
        spike_out_source199 = spike_out_source_array[199];
    end
    always @(spike_out_source_array[200]) begin 
        spike_out_source200 = spike_out_source_array[200];
    end
    always @(spike_out_source_array[201]) begin 
        spike_out_source201 = spike_out_source_array[201];
    end
    always @(spike_out_source_array[202]) begin 
        spike_out_source202 = spike_out_source_array[202];
    end
    always @(spike_out_source_array[203]) begin 
        spike_out_source203 = spike_out_source_array[203];
    end
    always @(spike_out_source_array[204]) begin 
        spike_out_source204 = spike_out_source_array[204];
    end
    always @(spike_out_source_array[205]) begin 
        spike_out_source205 = spike_out_source_array[205];
    end
    always @(spike_out_source_array[206]) begin 
        spike_out_source206 = spike_out_source_array[206];
    end
    always @(spike_out_source_array[207]) begin 
        spike_out_source207 = spike_out_source_array[207];
    end
    always @(spike_out_source_array[208]) begin 
        spike_out_source208 = spike_out_source_array[208];
    end
    always @(spike_out_source_array[209]) begin 
        spike_out_source209 = spike_out_source_array[209];
    end
    always @(spike_out_source_array[210]) begin 
        spike_out_source210 = spike_out_source_array[210];
    end
    always @(spike_out_source_array[211]) begin 
        spike_out_source211 = spike_out_source_array[211];
    end
    always @(spike_out_source_array[212]) begin 
        spike_out_source212 = spike_out_source_array[212];
    end
    always @(spike_out_source_array[213]) begin 
        spike_out_source213 = spike_out_source_array[213];
    end
    always @(spike_out_source_array[214]) begin 
        spike_out_source214 = spike_out_source_array[214];
    end
    always @(spike_out_source_array[215]) begin 
        spike_out_source215 = spike_out_source_array[215];
    end
    always @(spike_out_source_array[216]) begin 
        spike_out_source216 = spike_out_source_array[216];
    end
    always @(spike_out_source_array[217]) begin 
        spike_out_source217 = spike_out_source_array[217];
    end
    always @(spike_out_source_array[218]) begin 
        spike_out_source218 = spike_out_source_array[218];
    end
    always @(spike_out_source_array[219]) begin 
        spike_out_source219 = spike_out_source_array[219];
    end
    always @(spike_out_source_array[220]) begin 
        spike_out_source220 = spike_out_source_array[220];
    end
    always @(spike_out_source_array[221]) begin 
        spike_out_source221 = spike_out_source_array[221];
    end
    always @(spike_out_source_array[222]) begin 
        spike_out_source222 = spike_out_source_array[222];
    end
    always @(spike_out_source_array[223]) begin 
        spike_out_source223 = spike_out_source_array[223];
    end
    always @(spike_out_source_array[224]) begin 
        spike_out_source224 = spike_out_source_array[224];
    end
    always @(spike_out_source_array[225]) begin 
        spike_out_source225 = spike_out_source_array[225];
    end
    always @(spike_out_source_array[226]) begin 
        spike_out_source226 = spike_out_source_array[226];
    end
    always @(spike_out_source_array[227]) begin 
        spike_out_source227 = spike_out_source_array[227];
    end
    always @(spike_out_source_array[228]) begin 
        spike_out_source228 = spike_out_source_array[228];
    end
    always @(spike_out_source_array[229]) begin 
        spike_out_source229 = spike_out_source_array[229];
    end
    always @(spike_out_source_array[230]) begin 
        spike_out_source230 = spike_out_source_array[230];
    end
    always @(spike_out_source_array[231]) begin 
        spike_out_source231 = spike_out_source_array[231];
    end
    always @(spike_out_source_array[232]) begin 
        spike_out_source232 = spike_out_source_array[232];
    end
    always @(spike_out_source_array[233]) begin 
        spike_out_source233 = spike_out_source_array[233];
    end
    always @(spike_out_source_array[234]) begin 
        spike_out_source234 = spike_out_source_array[234];
    end
    always @(spike_out_source_array[235]) begin 
        spike_out_source235 = spike_out_source_array[235];
    end
    always @(spike_out_source_array[236]) begin 
        spike_out_source236 = spike_out_source_array[236];
    end
    always @(spike_out_source_array[237]) begin 
        spike_out_source237 = spike_out_source_array[237];
    end
    always @(spike_out_source_array[238]) begin 
        spike_out_source238 = spike_out_source_array[238];
    end
    always @(spike_out_source_array[239]) begin 
        spike_out_source239 = spike_out_source_array[239];
    end
    always @(spike_out_source_array[240]) begin 
        spike_out_source240 = spike_out_source_array[240];
    end
    always @(spike_out_source_array[241]) begin 
        spike_out_source241 = spike_out_source_array[241];
    end
    always @(spike_out_source_array[242]) begin 
        spike_out_source242 = spike_out_source_array[242];
    end
    always @(spike_out_source_array[243]) begin 
        spike_out_source243 = spike_out_source_array[243];
    end
    always @(spike_out_source_array[244]) begin 
        spike_out_source244 = spike_out_source_array[244];
    end
    always @(spike_out_source_array[245]) begin 
        spike_out_source245 = spike_out_source_array[245];
    end
    always @(spike_out_source_array[246]) begin 
        spike_out_source246 = spike_out_source_array[246];
    end
    always @(spike_out_source_array[247]) begin 
        spike_out_source247 = spike_out_source_array[247];
    end
    always @(spike_out_source_array[248]) begin 
        spike_out_source248 = spike_out_source_array[248];
    end
    always @(spike_out_source_array[249]) begin 
        spike_out_source249 = spike_out_source_array[249];
    end
    always @(spike_out_source_array[250]) begin 
        spike_out_source250 = spike_out_source_array[250];
    end
    always @(spike_out_source_array[251]) begin 
        spike_out_source251 = spike_out_source_array[251];
    end
    always @(spike_out_source_array[252]) begin 
        spike_out_source252 = spike_out_source_array[252];
    end
    always @(spike_out_source_array[253]) begin 
        spike_out_source253 = spike_out_source_array[253];
    end
    always @(spike_out_source_array[254]) begin 
        spike_out_source254 = spike_out_source_array[254];
    end
    always @(spike_out_source_array[255]) begin 
        spike_out_source255 = spike_out_source_array[255];
    end
    always @(spike_out_source_array[256]) begin 
        spike_out_source256 = spike_out_source_array[256];
    end
    always @(spike_out_source_array[257]) begin 
        spike_out_source257 = spike_out_source_array[257];
    end
    always @(spike_out_source_array[258]) begin 
        spike_out_source258 = spike_out_source_array[258];
    end
    always @(spike_out_source_array[259]) begin 
        spike_out_source259 = spike_out_source_array[259];
    end
    always @(spike_out_source_array[260]) begin 
        spike_out_source260 = spike_out_source_array[260];
    end
    always @(spike_out_source_array[261]) begin 
        spike_out_source261 = spike_out_source_array[261];
    end
    always @(spike_out_source_array[262]) begin 
        spike_out_source262 = spike_out_source_array[262];
    end
    always @(spike_out_source_array[263]) begin 
        spike_out_source263 = spike_out_source_array[263];
    end
    always @(spike_out_source_array[264]) begin 
        spike_out_source264 = spike_out_source_array[264];
    end
    always @(spike_out_source_array[265]) begin 
        spike_out_source265 = spike_out_source_array[265];
    end
    always @(spike_out_source_array[266]) begin 
        spike_out_source266 = spike_out_source_array[266];
    end
    always @(spike_out_source_array[267]) begin 
        spike_out_source267 = spike_out_source_array[267];
    end
    always @(spike_out_source_array[268]) begin 
        spike_out_source268 = spike_out_source_array[268];
    end
    always @(spike_out_source_array[269]) begin 
        spike_out_source269 = spike_out_source_array[269];
    end
    always @(spike_out_source_array[270]) begin 
        spike_out_source270 = spike_out_source_array[270];
    end
    always @(spike_out_source_array[271]) begin 
        spike_out_source271 = spike_out_source_array[271];
    end
    always @(spike_out_source_array[272]) begin 
        spike_out_source272 = spike_out_source_array[272];
    end
    always @(spike_out_source_array[273]) begin 
        spike_out_source273 = spike_out_source_array[273];
    end
    always @(spike_out_source_array[274]) begin 
        spike_out_source274 = spike_out_source_array[274];
    end
    always @(spike_out_source_array[275]) begin 
        spike_out_source275 = spike_out_source_array[275];
    end
    always @(spike_out_source_array[276]) begin 
        spike_out_source276 = spike_out_source_array[276];
    end
    always @(spike_out_source_array[277]) begin 
        spike_out_source277 = spike_out_source_array[277];
    end
    always @(spike_out_source_array[278]) begin 
        spike_out_source278 = spike_out_source_array[278];
    end
    always @(spike_out_source_array[279]) begin 
        spike_out_source279 = spike_out_source_array[279];
    end
    always @(spike_out_source_array[280]) begin 
        spike_out_source280 = spike_out_source_array[280];
    end
    always @(spike_out_source_array[281]) begin 
        spike_out_source281 = spike_out_source_array[281];
    end
    always @(spike_out_source_array[282]) begin 
        spike_out_source282 = spike_out_source_array[282];
    end
    always @(spike_out_source_array[283]) begin 
        spike_out_source283 = spike_out_source_array[283];
    end
    always @(spike_out_source_array[284]) begin 
        spike_out_source284 = spike_out_source_array[284];
    end
    always @(spike_out_source_array[285]) begin 
        spike_out_source285 = spike_out_source_array[285];
    end
    always @(spike_out_source_array[286]) begin 
        spike_out_source286 = spike_out_source_array[286];
    end
    always @(spike_out_source_array[287]) begin 
        spike_out_source287 = spike_out_source_array[287];
    end
    always @(spike_out_source_array[288]) begin 
        spike_out_source288 = spike_out_source_array[288];
    end
    always @(spike_out_source_array[289]) begin 
        spike_out_source289 = spike_out_source_array[289];
    end
    always @(spike_out_source_array[290]) begin 
        spike_out_source290 = spike_out_source_array[290];
    end
    always @(spike_out_source_array[291]) begin 
        spike_out_source291 = spike_out_source_array[291];
    end
    always @(spike_out_source_array[292]) begin 
        spike_out_source292 = spike_out_source_array[292];
    end
    always @(spike_out_source_array[293]) begin 
        spike_out_source293 = spike_out_source_array[293];
    end
    always @(spike_out_source_array[294]) begin 
        spike_out_source294 = spike_out_source_array[294];
    end
    always @(spike_out_source_array[295]) begin 
        spike_out_source295 = spike_out_source_array[295];
    end
    always @(spike_out_source_array[296]) begin 
        spike_out_source296 = spike_out_source_array[296];
    end
    always @(spike_out_source_array[297]) begin 
        spike_out_source297 = spike_out_source_array[297];
    end
    always @(spike_out_source_array[298]) begin 
        spike_out_source298 = spike_out_source_array[298];
    end
    always @(spike_out_source_array[299]) begin 
        spike_out_source299 = spike_out_source_array[299];
    end
    always @(spike_out_source_array[300]) begin 
        spike_out_source300 = spike_out_source_array[300];
    end
    always @(spike_out_source_array[301]) begin 
        spike_out_source301 = spike_out_source_array[301];
    end
    always @(spike_out_source_array[302]) begin 
        spike_out_source302 = spike_out_source_array[302];
    end
    always @(spike_out_source_array[303]) begin 
        spike_out_source303 = spike_out_source_array[303];
    end
    always @(spike_out_source_array[304]) begin 
        spike_out_source304 = spike_out_source_array[304];
    end
    always @(spike_out_source_array[305]) begin 
        spike_out_source305 = spike_out_source_array[305];
    end
    always @(spike_out_source_array[306]) begin 
        spike_out_source306 = spike_out_source_array[306];
    end
    always @(spike_out_source_array[307]) begin 
        spike_out_source307 = spike_out_source_array[307];
    end
    always @(spike_out_source_array[308]) begin 
        spike_out_source308 = spike_out_source_array[308];
    end
    always @(spike_out_source_array[309]) begin 
        spike_out_source309 = spike_out_source_array[309];
    end
    always @(spike_out_source_array[310]) begin 
        spike_out_source310 = spike_out_source_array[310];
    end
    always @(spike_out_source_array[311]) begin 
        spike_out_source311 = spike_out_source_array[311];
    end
    always @(spike_out_source_array[312]) begin 
        spike_out_source312 = spike_out_source_array[312];
    end
    always @(spike_out_source_array[313]) begin 
        spike_out_source313 = spike_out_source_array[313];
    end
    always @(spike_out_source_array[314]) begin 
        spike_out_source314 = spike_out_source_array[314];
    end
    always @(spike_out_source_array[315]) begin 
        spike_out_source315 = spike_out_source_array[315];
    end
    always @(spike_out_source_array[316]) begin 
        spike_out_source316 = spike_out_source_array[316];
    end
    always @(spike_out_source_array[317]) begin 
        spike_out_source317 = spike_out_source_array[317];
    end
    always @(spike_out_source_array[318]) begin 
        spike_out_source318 = spike_out_source_array[318];
    end
    always @(spike_out_source_array[319]) begin 
        spike_out_source319 = spike_out_source_array[319];
    end
    always @(spike_out_source_array[320]) begin 
        spike_out_source320 = spike_out_source_array[320];
    end
    always @(spike_out_source_array[321]) begin 
        spike_out_source321 = spike_out_source_array[321];
    end
    always @(spike_out_source_array[322]) begin 
        spike_out_source322 = spike_out_source_array[322];
    end
    always @(spike_out_source_array[323]) begin 
        spike_out_source323 = spike_out_source_array[323];
    end
    always @(spike_out_source_array[324]) begin 
        spike_out_source324 = spike_out_source_array[324];
    end
    always @(spike_out_source_array[325]) begin 
        spike_out_source325 = spike_out_source_array[325];
    end
    always @(spike_out_source_array[326]) begin 
        spike_out_source326 = spike_out_source_array[326];
    end
    always @(spike_out_source_array[327]) begin 
        spike_out_source327 = spike_out_source_array[327];
    end
    always @(spike_out_source_array[328]) begin 
        spike_out_source328 = spike_out_source_array[328];
    end
    always @(spike_out_source_array[329]) begin 
        spike_out_source329 = spike_out_source_array[329];
    end
    always @(spike_out_source_array[330]) begin 
        spike_out_source330 = spike_out_source_array[330];
    end
    always @(spike_out_source_array[331]) begin 
        spike_out_source331 = spike_out_source_array[331];
    end
    always @(spike_out_source_array[332]) begin 
        spike_out_source332 = spike_out_source_array[332];
    end
    always @(spike_out_source_array[333]) begin 
        spike_out_source333 = spike_out_source_array[333];
    end
    always @(spike_out_source_array[334]) begin 
        spike_out_source334 = spike_out_source_array[334];
    end
    always @(spike_out_source_array[335]) begin 
        spike_out_source335 = spike_out_source_array[335];
    end
    always @(spike_out_source_array[336]) begin 
        spike_out_source336 = spike_out_source_array[336];
    end
    always @(spike_out_source_array[337]) begin 
        spike_out_source337 = spike_out_source_array[337];
    end
    always @(spike_out_source_array[338]) begin 
        spike_out_source338 = spike_out_source_array[338];
    end
    always @(spike_out_source_array[339]) begin 
        spike_out_source339 = spike_out_source_array[339];
    end
    always @(spike_out_source_array[340]) begin 
        spike_out_source340 = spike_out_source_array[340];
    end
    always @(spike_out_source_array[341]) begin 
        spike_out_source341 = spike_out_source_array[341];
    end
    always @(spike_out_source_array[342]) begin 
        spike_out_source342 = spike_out_source_array[342];
    end
    always @(spike_out_source_array[343]) begin 
        spike_out_source343 = spike_out_source_array[343];
    end
    always @(spike_out_source_array[344]) begin 
        spike_out_source344 = spike_out_source_array[344];
    end
    always @(spike_out_source_array[345]) begin 
        spike_out_source345 = spike_out_source_array[345];
    end
    always @(spike_out_source_array[346]) begin 
        spike_out_source346 = spike_out_source_array[346];
    end
    always @(spike_out_source_array[347]) begin 
        spike_out_source347 = spike_out_source_array[347];
    end
    always @(spike_out_source_array[348]) begin 
        spike_out_source348 = spike_out_source_array[348];
    end
    always @(spike_out_source_array[349]) begin 
        spike_out_source349 = spike_out_source_array[349];
    end
    always @(spike_out_source_array[350]) begin 
        spike_out_source350 = spike_out_source_array[350];
    end
    always @(spike_out_source_array[351]) begin 
        spike_out_source351 = spike_out_source_array[351];
    end
    always @(spike_out_source_array[352]) begin 
        spike_out_source352 = spike_out_source_array[352];
    end
    always @(spike_out_source_array[353]) begin 
        spike_out_source353 = spike_out_source_array[353];
    end
    always @(spike_out_source_array[354]) begin 
        spike_out_source354 = spike_out_source_array[354];
    end
    always @(spike_out_source_array[355]) begin 
        spike_out_source355 = spike_out_source_array[355];
    end
    always @(spike_out_source_array[356]) begin 
        spike_out_source356 = spike_out_source_array[356];
    end
    always @(spike_out_source_array[357]) begin 
        spike_out_source357 = spike_out_source_array[357];
    end
    always @(spike_out_source_array[358]) begin 
        spike_out_source358 = spike_out_source_array[358];
    end
    always @(spike_out_source_array[359]) begin 
        spike_out_source359 = spike_out_source_array[359];
    end
    always @(spike_out_source_array[360]) begin 
        spike_out_source360 = spike_out_source_array[360];
    end
    always @(spike_out_source_array[361]) begin 
        spike_out_source361 = spike_out_source_array[361];
    end
    always @(spike_out_source_array[362]) begin 
        spike_out_source362 = spike_out_source_array[362];
    end
    always @(spike_out_source_array[363]) begin 
        spike_out_source363 = spike_out_source_array[363];
    end
    always @(spike_out_source_array[364]) begin 
        spike_out_source364 = spike_out_source_array[364];
    end
    always @(spike_out_source_array[365]) begin 
        spike_out_source365 = spike_out_source_array[365];
    end
    always @(spike_out_source_array[366]) begin 
        spike_out_source366 = spike_out_source_array[366];
    end
    always @(spike_out_source_array[367]) begin 
        spike_out_source367 = spike_out_source_array[367];
    end
    always @(spike_out_source_array[368]) begin 
        spike_out_source368 = spike_out_source_array[368];
    end
    always @(spike_out_source_array[369]) begin 
        spike_out_source369 = spike_out_source_array[369];
    end
    always @(spike_out_source_array[370]) begin 
        spike_out_source370 = spike_out_source_array[370];
    end
    always @(spike_out_source_array[371]) begin 
        spike_out_source371 = spike_out_source_array[371];
    end
    always @(spike_out_source_array[372]) begin 
        spike_out_source372 = spike_out_source_array[372];
    end
    always @(spike_out_source_array[373]) begin 
        spike_out_source373 = spike_out_source_array[373];
    end
    always @(spike_out_source_array[374]) begin 
        spike_out_source374 = spike_out_source_array[374];
    end
    always @(spike_out_source_array[375]) begin 
        spike_out_source375 = spike_out_source_array[375];
    end
    always @(spike_out_source_array[376]) begin 
        spike_out_source376 = spike_out_source_array[376];
    end
    always @(spike_out_source_array[377]) begin 
        spike_out_source377 = spike_out_source_array[377];
    end
    always @(spike_out_source_array[378]) begin 
        spike_out_source378 = spike_out_source_array[378];
    end
    always @(spike_out_source_array[379]) begin 
        spike_out_source379 = spike_out_source_array[379];
    end
    always @(spike_out_source_array[380]) begin 
        spike_out_source380 = spike_out_source_array[380];
    end
    always @(spike_out_source_array[381]) begin 
        spike_out_source381 = spike_out_source_array[381];
    end
    always @(spike_out_source_array[382]) begin 
        spike_out_source382 = spike_out_source_array[382];
    end
    always @(spike_out_source_array[383]) begin 
        spike_out_source383 = spike_out_source_array[383];
    end
    always @(spike_out_source_array[384]) begin 
        spike_out_source384 = spike_out_source_array[384];
    end
    always @(spike_out_source_array[385]) begin 
        spike_out_source385 = spike_out_source_array[385];
    end
    always @(spike_out_source_array[386]) begin 
        spike_out_source386 = spike_out_source_array[386];
    end
    always @(spike_out_source_array[387]) begin 
        spike_out_source387 = spike_out_source_array[387];
    end
    always @(spike_out_source_array[388]) begin 
        spike_out_source388 = spike_out_source_array[388];
    end
    always @(spike_out_source_array[389]) begin 
        spike_out_source389 = spike_out_source_array[389];
    end
    always @(spike_out_source_array[390]) begin 
        spike_out_source390 = spike_out_source_array[390];
    end
    always @(spike_out_source_array[391]) begin 
        spike_out_source391 = spike_out_source_array[391];
    end
    always @(spike_out_source_array[392]) begin 
        spike_out_source392 = spike_out_source_array[392];
    end
    always @(spike_out_source_array[393]) begin 
        spike_out_source393 = spike_out_source_array[393];
    end
    always @(spike_out_source_array[394]) begin 
        spike_out_source394 = spike_out_source_array[394];
    end
    always @(spike_out_source_array[395]) begin 
        spike_out_source395 = spike_out_source_array[395];
    end
    always @(spike_out_source_array[396]) begin 
        spike_out_source396 = spike_out_source_array[396];
    end
    always @(spike_out_source_array[397]) begin 
        spike_out_source397 = spike_out_source_array[397];
    end
    always @(spike_out_source_array[398]) begin 
        spike_out_source398 = spike_out_source_array[398];
    end
    always @(spike_out_source_array[399]) begin 
        spike_out_source399 = spike_out_source_array[399];
    end
    always @(spike_out_source_array[400]) begin 
        spike_out_source400 = spike_out_source_array[400];
    end
    always @(spike_out_source_array[401]) begin 
        spike_out_source401 = spike_out_source_array[401];
    end
    always @(spike_out_source_array[402]) begin 
        spike_out_source402 = spike_out_source_array[402];
    end
    always @(spike_out_source_array[403]) begin 
        spike_out_source403 = spike_out_source_array[403];
    end
    always @(spike_out_source_array[404]) begin 
        spike_out_source404 = spike_out_source_array[404];
    end
    always @(spike_out_source_array[405]) begin 
        spike_out_source405 = spike_out_source_array[405];
    end
    always @(spike_out_source_array[406]) begin 
        spike_out_source406 = spike_out_source_array[406];
    end
    always @(spike_out_source_array[407]) begin 
        spike_out_source407 = spike_out_source_array[407];
    end
    always @(spike_out_source_array[408]) begin 
        spike_out_source408 = spike_out_source_array[408];
    end
    always @(spike_out_source_array[409]) begin 
        spike_out_source409 = spike_out_source_array[409];
    end
    always @(spike_out_source_array[410]) begin 
        spike_out_source410 = spike_out_source_array[410];
    end
    always @(spike_out_source_array[411]) begin 
        spike_out_source411 = spike_out_source_array[411];
    end
    always @(spike_out_source_array[412]) begin 
        spike_out_source412 = spike_out_source_array[412];
    end
    always @(spike_out_source_array[413]) begin 
        spike_out_source413 = spike_out_source_array[413];
    end
    always @(spike_out_source_array[414]) begin 
        spike_out_source414 = spike_out_source_array[414];
    end
    always @(spike_out_source_array[415]) begin 
        spike_out_source415 = spike_out_source_array[415];
    end
    always @(spike_out_source_array[416]) begin 
        spike_out_source416 = spike_out_source_array[416];
    end
    always @(spike_out_source_array[417]) begin 
        spike_out_source417 = spike_out_source_array[417];
    end
    always @(spike_out_source_array[418]) begin 
        spike_out_source418 = spike_out_source_array[418];
    end
    always @(spike_out_source_array[419]) begin 
        spike_out_source419 = spike_out_source_array[419];
    end
    always @(spike_out_source_array[420]) begin 
        spike_out_source420 = spike_out_source_array[420];
    end
    always @(spike_out_source_array[421]) begin 
        spike_out_source421 = spike_out_source_array[421];
    end
    always @(spike_out_source_array[422]) begin 
        spike_out_source422 = spike_out_source_array[422];
    end
    always @(spike_out_source_array[423]) begin 
        spike_out_source423 = spike_out_source_array[423];
    end
    always @(spike_out_source_array[424]) begin 
        spike_out_source424 = spike_out_source_array[424];
    end
    always @(spike_out_source_array[425]) begin 
        spike_out_source425 = spike_out_source_array[425];
    end
    always @(spike_out_source_array[426]) begin 
        spike_out_source426 = spike_out_source_array[426];
    end
    always @(spike_out_source_array[427]) begin 
        spike_out_source427 = spike_out_source_array[427];
    end
    always @(spike_out_source_array[428]) begin 
        spike_out_source428 = spike_out_source_array[428];
    end
    always @(spike_out_source_array[429]) begin 
        spike_out_source429 = spike_out_source_array[429];
    end
    always @(spike_out_source_array[430]) begin 
        spike_out_source430 = spike_out_source_array[430];
    end
    always @(spike_out_source_array[431]) begin 
        spike_out_source431 = spike_out_source_array[431];
    end
    always @(spike_out_source_array[432]) begin 
        spike_out_source432 = spike_out_source_array[432];
    end
    always @(spike_out_source_array[433]) begin 
        spike_out_source433 = spike_out_source_array[433];
    end
    always @(spike_out_source_array[434]) begin 
        spike_out_source434 = spike_out_source_array[434];
    end
    always @(spike_out_source_array[435]) begin 
        spike_out_source435 = spike_out_source_array[435];
    end
    always @(spike_out_source_array[436]) begin 
        spike_out_source436 = spike_out_source_array[436];
    end
    always @(spike_out_source_array[437]) begin 
        spike_out_source437 = spike_out_source_array[437];
    end
    always @(spike_out_source_array[438]) begin 
        spike_out_source438 = spike_out_source_array[438];
    end
    always @(spike_out_source_array[439]) begin 
        spike_out_source439 = spike_out_source_array[439];
    end
    always @(spike_out_source_array[440]) begin 
        spike_out_source440 = spike_out_source_array[440];
    end
    always @(spike_out_source_array[441]) begin 
        spike_out_source441 = spike_out_source_array[441];
    end
    always @(spike_out_source_array[442]) begin 
        spike_out_source442 = spike_out_source_array[442];
    end
    always @(spike_out_source_array[443]) begin 
        spike_out_source443 = spike_out_source_array[443];
    end
    always @(spike_out_source_array[444]) begin 
        spike_out_source444 = spike_out_source_array[444];
    end
    always @(spike_out_source_array[445]) begin 
        spike_out_source445 = spike_out_source_array[445];
    end
    always @(spike_out_source_array[446]) begin 
        spike_out_source446 = spike_out_source_array[446];
    end
    always @(spike_out_source_array[447]) begin 
        spike_out_source447 = spike_out_source_array[447];
    end
    always @(spike_out_source_array[448]) begin 
        spike_out_source448 = spike_out_source_array[448];
    end
    always @(spike_out_source_array[449]) begin 
        spike_out_source449 = spike_out_source_array[449];
    end
    always @(spike_out_source_array[450]) begin 
        spike_out_source450 = spike_out_source_array[450];
    end
    always @(spike_out_source_array[451]) begin 
        spike_out_source451 = spike_out_source_array[451];
    end
    always @(spike_out_source_array[452]) begin 
        spike_out_source452 = spike_out_source_array[452];
    end
    always @(spike_out_source_array[453]) begin 
        spike_out_source453 = spike_out_source_array[453];
    end
    always @(spike_out_source_array[454]) begin 
        spike_out_source454 = spike_out_source_array[454];
    end
    always @(spike_out_source_array[455]) begin 
        spike_out_source455 = spike_out_source_array[455];
    end
    always @(spike_out_source_array[456]) begin 
        spike_out_source456 = spike_out_source_array[456];
    end
    always @(spike_out_source_array[457]) begin 
        spike_out_source457 = spike_out_source_array[457];
    end
    always @(spike_out_source_array[458]) begin 
        spike_out_source458 = spike_out_source_array[458];
    end
    always @(spike_out_source_array[459]) begin 
        spike_out_source459 = spike_out_source_array[459];
    end
    always @(spike_out_source_array[460]) begin 
        spike_out_source460 = spike_out_source_array[460];
    end
    always @(spike_out_source_array[461]) begin 
        spike_out_source461 = spike_out_source_array[461];
    end
    always @(spike_out_source_array[462]) begin 
        spike_out_source462 = spike_out_source_array[462];
    end
    always @(spike_out_source_array[463]) begin 
        spike_out_source463 = spike_out_source_array[463];
    end
    always @(spike_out_source_array[464]) begin 
        spike_out_source464 = spike_out_source_array[464];
    end
    always @(spike_out_source_array[465]) begin 
        spike_out_source465 = spike_out_source_array[465];
    end
    always @(spike_out_source_array[466]) begin 
        spike_out_source466 = spike_out_source_array[466];
    end
    always @(spike_out_source_array[467]) begin 
        spike_out_source467 = spike_out_source_array[467];
    end
    always @(spike_out_source_array[468]) begin 
        spike_out_source468 = spike_out_source_array[468];
    end
    always @(spike_out_source_array[469]) begin 
        spike_out_source469 = spike_out_source_array[469];
    end
    always @(spike_out_source_array[470]) begin 
        spike_out_source470 = spike_out_source_array[470];
    end
    always @(spike_out_source_array[471]) begin 
        spike_out_source471 = spike_out_source_array[471];
    end
    always @(spike_out_source_array[472]) begin 
        spike_out_source472 = spike_out_source_array[472];
    end
    always @(spike_out_source_array[473]) begin 
        spike_out_source473 = spike_out_source_array[473];
    end
    always @(spike_out_source_array[474]) begin 
        spike_out_source474 = spike_out_source_array[474];
    end
    always @(spike_out_source_array[475]) begin 
        spike_out_source475 = spike_out_source_array[475];
    end
    always @(spike_out_source_array[476]) begin 
        spike_out_source476 = spike_out_source_array[476];
    end
    always @(spike_out_source_array[477]) begin 
        spike_out_source477 = spike_out_source_array[477];
    end
    always @(spike_out_source_array[478]) begin 
        spike_out_source478 = spike_out_source_array[478];
    end
    always @(spike_out_source_array[479]) begin 
        spike_out_source479 = spike_out_source_array[479];
    end
    always @(spike_out_source_array[480]) begin 
        spike_out_source480 = spike_out_source_array[480];
    end
    always @(spike_out_source_array[481]) begin 
        spike_out_source481 = spike_out_source_array[481];
    end
    always @(spike_out_source_array[482]) begin 
        spike_out_source482 = spike_out_source_array[482];
    end
    always @(spike_out_source_array[483]) begin 
        spike_out_source483 = spike_out_source_array[483];
    end
    always @(spike_out_source_array[484]) begin 
        spike_out_source484 = spike_out_source_array[484];
    end
    always @(spike_out_source_array[485]) begin 
        spike_out_source485 = spike_out_source_array[485];
    end
    always @(spike_out_source_array[486]) begin 
        spike_out_source486 = spike_out_source_array[486];
    end
    always @(spike_out_source_array[487]) begin 
        spike_out_source487 = spike_out_source_array[487];
    end
    always @(spike_out_source_array[488]) begin 
        spike_out_source488 = spike_out_source_array[488];
    end
    always @(spike_out_source_array[489]) begin 
        spike_out_source489 = spike_out_source_array[489];
    end
    always @(spike_out_source_array[490]) begin 
        spike_out_source490 = spike_out_source_array[490];
    end
    always @(spike_out_source_array[491]) begin 
        spike_out_source491 = spike_out_source_array[491];
    end
    always @(spike_out_source_array[492]) begin 
        spike_out_source492 = spike_out_source_array[492];
    end
    always @(spike_out_source_array[493]) begin 
        spike_out_source493 = spike_out_source_array[493];
    end
    always @(spike_out_source_array[494]) begin 
        spike_out_source494 = spike_out_source_array[494];
    end
    always @(spike_out_source_array[495]) begin 
        spike_out_source495 = spike_out_source_array[495];
    end
    always @(spike_out_source_array[496]) begin 
        spike_out_source496 = spike_out_source_array[496];
    end
    always @(spike_out_source_array[497]) begin 
        spike_out_source497 = spike_out_source_array[497];
    end
    always @(spike_out_source_array[498]) begin 
        spike_out_source498 = spike_out_source_array[498];
    end
    always @(spike_out_source_array[499]) begin 
        spike_out_source499 = spike_out_source_array[499];
    end
    always @(spike_out_source_array[500]) begin 
        spike_out_source500 = spike_out_source_array[500];
    end
    always @(spike_out_source_array[501]) begin 
        spike_out_source501 = spike_out_source_array[501];
    end
    always @(spike_out_source_array[502]) begin 
        spike_out_source502 = spike_out_source_array[502];
    end
    always @(spike_out_source_array[503]) begin 
        spike_out_source503 = spike_out_source_array[503];
    end
    always @(spike_out_source_array[504]) begin 
        spike_out_source504 = spike_out_source_array[504];
    end
    always @(spike_out_source_array[505]) begin 
        spike_out_source505 = spike_out_source_array[505];
    end
    always @(spike_out_source_array[506]) begin 
        spike_out_source506 = spike_out_source_array[506];
    end
    always @(spike_out_source_array[507]) begin 
        spike_out_source507 = spike_out_source_array[507];
    end
    always @(spike_out_source_array[508]) begin 
        spike_out_source508 = spike_out_source_array[508];
    end
    always @(spike_out_source_array[509]) begin 
        spike_out_source509 = spike_out_source_array[509];
    end
    always @(spike_out_source_array[510]) begin 
        spike_out_source510 = spike_out_source_array[510];
    end
    always @(spike_out_source_array[511]) begin 
        spike_out_source511 = spike_out_source_array[511];
    end
    always @(spike_out_source_array[512]) begin 
        spike_out_source512 = spike_out_source_array[512];
    end
    always @(spike_out_source_array[513]) begin 
        spike_out_source513 = spike_out_source_array[513];
    end
    always @(spike_out_source_array[514]) begin 
        spike_out_source514 = spike_out_source_array[514];
    end
    always @(spike_out_source_array[515]) begin 
        spike_out_source515 = spike_out_source_array[515];
    end
    always @(spike_out_source_array[516]) begin 
        spike_out_source516 = spike_out_source_array[516];
    end
    always @(spike_out_source_array[517]) begin 
        spike_out_source517 = spike_out_source_array[517];
    end
    always @(spike_out_source_array[518]) begin 
        spike_out_source518 = spike_out_source_array[518];
    end
    always @(spike_out_source_array[519]) begin 
        spike_out_source519 = spike_out_source_array[519];
    end
    always @(spike_out_source_array[520]) begin 
        spike_out_source520 = spike_out_source_array[520];
    end
    always @(spike_out_source_array[521]) begin 
        spike_out_source521 = spike_out_source_array[521];
    end
    always @(spike_out_source_array[522]) begin 
        spike_out_source522 = spike_out_source_array[522];
    end
    always @(spike_out_source_array[523]) begin 
        spike_out_source523 = spike_out_source_array[523];
    end
    always @(spike_out_source_array[524]) begin 
        spike_out_source524 = spike_out_source_array[524];
    end
    always @(spike_out_source_array[525]) begin 
        spike_out_source525 = spike_out_source_array[525];
    end
    always @(spike_out_source_array[526]) begin 
        spike_out_source526 = spike_out_source_array[526];
    end
    always @(spike_out_source_array[527]) begin 
        spike_out_source527 = spike_out_source_array[527];
    end
    always @(spike_out_source_array[528]) begin 
        spike_out_source528 = spike_out_source_array[528];
    end
    always @(spike_out_source_array[529]) begin 
        spike_out_source529 = spike_out_source_array[529];
    end
    always @(spike_out_source_array[530]) begin 
        spike_out_source530 = spike_out_source_array[530];
    end
    always @(spike_out_source_array[531]) begin 
        spike_out_source531 = spike_out_source_array[531];
    end
    always @(spike_out_source_array[532]) begin 
        spike_out_source532 = spike_out_source_array[532];
    end
    always @(spike_out_source_array[533]) begin 
        spike_out_source533 = spike_out_source_array[533];
    end
    always @(spike_out_source_array[534]) begin 
        spike_out_source534 = spike_out_source_array[534];
    end
    always @(spike_out_source_array[535]) begin 
        spike_out_source535 = spike_out_source_array[535];
    end
    always @(spike_out_source_array[536]) begin 
        spike_out_source536 = spike_out_source_array[536];
    end
    always @(spike_out_source_array[537]) begin 
        spike_out_source537 = spike_out_source_array[537];
    end
    always @(spike_out_source_array[538]) begin 
        spike_out_source538 = spike_out_source_array[538];
    end
    always @(spike_out_source_array[539]) begin 
        spike_out_source539 = spike_out_source_array[539];
    end
    always @(spike_out_source_array[540]) begin 
        spike_out_source540 = spike_out_source_array[540];
    end
    always @(spike_out_source_array[541]) begin 
        spike_out_source541 = spike_out_source_array[541];
    end
    always @(spike_out_source_array[542]) begin 
        spike_out_source542 = spike_out_source_array[542];
    end
    always @(spike_out_source_array[543]) begin 
        spike_out_source543 = spike_out_source_array[543];
    end
    always @(spike_out_source_array[544]) begin 
        spike_out_source544 = spike_out_source_array[544];
    end
    always @(spike_out_source_array[545]) begin 
        spike_out_source545 = spike_out_source_array[545];
    end
    always @(spike_out_source_array[546]) begin 
        spike_out_source546 = spike_out_source_array[546];
    end
    always @(spike_out_source_array[547]) begin 
        spike_out_source547 = spike_out_source_array[547];
    end
    always @(spike_out_source_array[548]) begin 
        spike_out_source548 = spike_out_source_array[548];
    end
    always @(spike_out_source_array[549]) begin 
        spike_out_source549 = spike_out_source_array[549];
    end
    always @(spike_out_source_array[550]) begin 
        spike_out_source550 = spike_out_source_array[550];
    end
    always @(spike_out_source_array[551]) begin 
        spike_out_source551 = spike_out_source_array[551];
    end
    always @(spike_out_source_array[552]) begin 
        spike_out_source552 = spike_out_source_array[552];
    end
    always @(spike_out_source_array[553]) begin 
        spike_out_source553 = spike_out_source_array[553];
    end
    always @(spike_out_source_array[554]) begin 
        spike_out_source554 = spike_out_source_array[554];
    end
    always @(spike_out_source_array[555]) begin 
        spike_out_source555 = spike_out_source_array[555];
    end
    always @(spike_out_source_array[556]) begin 
        spike_out_source556 = spike_out_source_array[556];
    end
    always @(spike_out_source_array[557]) begin 
        spike_out_source557 = spike_out_source_array[557];
    end
    always @(spike_out_source_array[558]) begin 
        spike_out_source558 = spike_out_source_array[558];
    end
    always @(spike_out_source_array[559]) begin 
        spike_out_source559 = spike_out_source_array[559];
    end
    always @(spike_out_source_array[560]) begin 
        spike_out_source560 = spike_out_source_array[560];
    end
    always @(spike_out_source_array[561]) begin 
        spike_out_source561 = spike_out_source_array[561];
    end
    always @(spike_out_source_array[562]) begin 
        spike_out_source562 = spike_out_source_array[562];
    end
    always @(spike_out_source_array[563]) begin 
        spike_out_source563 = spike_out_source_array[563];
    end
    always @(spike_out_source_array[564]) begin 
        spike_out_source564 = spike_out_source_array[564];
    end
    always @(spike_out_source_array[565]) begin 
        spike_out_source565 = spike_out_source_array[565];
    end
    always @(spike_out_source_array[566]) begin 
        spike_out_source566 = spike_out_source_array[566];
    end
    always @(spike_out_source_array[567]) begin 
        spike_out_source567 = spike_out_source_array[567];
    end
    always @(spike_out_source_array[568]) begin 
        spike_out_source568 = spike_out_source_array[568];
    end
    always @(spike_out_source_array[569]) begin 
        spike_out_source569 = spike_out_source_array[569];
    end
    always @(spike_out_source_array[570]) begin 
        spike_out_source570 = spike_out_source_array[570];
    end
    always @(spike_out_source_array[571]) begin 
        spike_out_source571 = spike_out_source_array[571];
    end
    always @(spike_out_source_array[572]) begin 
        spike_out_source572 = spike_out_source_array[572];
    end
    always @(spike_out_source_array[573]) begin 
        spike_out_source573 = spike_out_source_array[573];
    end
    always @(spike_out_source_array[574]) begin 
        spike_out_source574 = spike_out_source_array[574];
    end
    always @(spike_out_source_array[575]) begin 
        spike_out_source575 = spike_out_source_array[575];
    end
    always @(spike_out_source_array[576]) begin 
        spike_out_source576 = spike_out_source_array[576];
    end
    always @(spike_out_source_array[577]) begin 
        spike_out_source577 = spike_out_source_array[577];
    end
    always @(spike_out_source_array[578]) begin 
        spike_out_source578 = spike_out_source_array[578];
    end
    always @(spike_out_source_array[579]) begin 
        spike_out_source579 = spike_out_source_array[579];
    end
    always @(spike_out_source_array[580]) begin 
        spike_out_source580 = spike_out_source_array[580];
    end
    always @(spike_out_source_array[581]) begin 
        spike_out_source581 = spike_out_source_array[581];
    end
    always @(spike_out_source_array[582]) begin 
        spike_out_source582 = spike_out_source_array[582];
    end
    always @(spike_out_source_array[583]) begin 
        spike_out_source583 = spike_out_source_array[583];
    end
    always @(spike_out_source_array[584]) begin 
        spike_out_source584 = spike_out_source_array[584];
    end
    always @(spike_out_source_array[585]) begin 
        spike_out_source585 = spike_out_source_array[585];
    end
    always @(spike_out_source_array[586]) begin 
        spike_out_source586 = spike_out_source_array[586];
    end
    always @(spike_out_source_array[587]) begin 
        spike_out_source587 = spike_out_source_array[587];
    end
    always @(spike_out_source_array[588]) begin 
        spike_out_source588 = spike_out_source_array[588];
    end
    always @(spike_out_source_array[589]) begin 
        spike_out_source589 = spike_out_source_array[589];
    end
    always @(spike_out_source_array[590]) begin 
        spike_out_source590 = spike_out_source_array[590];
    end
    always @(spike_out_source_array[591]) begin 
        spike_out_source591 = spike_out_source_array[591];
    end
    always @(spike_out_source_array[592]) begin 
        spike_out_source592 = spike_out_source_array[592];
    end
    always @(spike_out_source_array[593]) begin 
        spike_out_source593 = spike_out_source_array[593];
    end
    always @(spike_out_source_array[594]) begin 
        spike_out_source594 = spike_out_source_array[594];
    end
    always @(spike_out_source_array[595]) begin 
        spike_out_source595 = spike_out_source_array[595];
    end
    always @(spike_out_source_array[596]) begin 
        spike_out_source596 = spike_out_source_array[596];
    end
    always @(spike_out_source_array[597]) begin 
        spike_out_source597 = spike_out_source_array[597];
    end
    always @(spike_out_source_array[598]) begin 
        spike_out_source598 = spike_out_source_array[598];
    end
    always @(spike_out_source_array[599]) begin 
        spike_out_source599 = spike_out_source_array[599];
    end
    always @(spike_out_source_array[600]) begin 
        spike_out_source600 = spike_out_source_array[600];
    end
    always @(spike_out_source_array[601]) begin 
        spike_out_source601 = spike_out_source_array[601];
    end
    always @(spike_out_source_array[602]) begin 
        spike_out_source602 = spike_out_source_array[602];
    end
    always @(spike_out_source_array[603]) begin 
        spike_out_source603 = spike_out_source_array[603];
    end
    always @(spike_out_source_array[604]) begin 
        spike_out_source604 = spike_out_source_array[604];
    end
    always @(spike_out_source_array[605]) begin 
        spike_out_source605 = spike_out_source_array[605];
    end
    always @(spike_out_source_array[606]) begin 
        spike_out_source606 = spike_out_source_array[606];
    end
    always @(spike_out_source_array[607]) begin 
        spike_out_source607 = spike_out_source_array[607];
    end
    always @(spike_out_source_array[608]) begin 
        spike_out_source608 = spike_out_source_array[608];
    end
    always @(spike_out_source_array[609]) begin 
        spike_out_source609 = spike_out_source_array[609];
    end
    always @(spike_out_source_array[610]) begin 
        spike_out_source610 = spike_out_source_array[610];
    end
    always @(spike_out_source_array[611]) begin 
        spike_out_source611 = spike_out_source_array[611];
    end
    always @(spike_out_source_array[612]) begin 
        spike_out_source612 = spike_out_source_array[612];
    end
    always @(spike_out_source_array[613]) begin 
        spike_out_source613 = spike_out_source_array[613];
    end
    always @(spike_out_source_array[614]) begin 
        spike_out_source614 = spike_out_source_array[614];
    end
    always @(spike_out_source_array[615]) begin 
        spike_out_source615 = spike_out_source_array[615];
    end
    always @(spike_out_source_array[616]) begin 
        spike_out_source616 = spike_out_source_array[616];
    end
    always @(spike_out_source_array[617]) begin 
        spike_out_source617 = spike_out_source_array[617];
    end
    always @(spike_out_source_array[618]) begin 
        spike_out_source618 = spike_out_source_array[618];
    end
    always @(spike_out_source_array[619]) begin 
        spike_out_source619 = spike_out_source_array[619];
    end
    always @(spike_out_source_array[620]) begin 
        spike_out_source620 = spike_out_source_array[620];
    end
    always @(spike_out_source_array[621]) begin 
        spike_out_source621 = spike_out_source_array[621];
    end
    always @(spike_out_source_array[622]) begin 
        spike_out_source622 = spike_out_source_array[622];
    end
    always @(spike_out_source_array[623]) begin 
        spike_out_source623 = spike_out_source_array[623];
    end
    always @(spike_out_source_array[624]) begin 
        spike_out_source624 = spike_out_source_array[624];
    end
    always @(spike_out_source_array[625]) begin 
        spike_out_source625 = spike_out_source_array[625];
    end
    always @(spike_out_source_array[626]) begin 
        spike_out_source626 = spike_out_source_array[626];
    end
    always @(spike_out_source_array[627]) begin 
        spike_out_source627 = spike_out_source_array[627];
    end
    always @(spike_out_source_array[628]) begin 
        spike_out_source628 = spike_out_source_array[628];
    end
    always @(spike_out_source_array[629]) begin 
        spike_out_source629 = spike_out_source_array[629];
    end
    always @(spike_out_source_array[630]) begin 
        spike_out_source630 = spike_out_source_array[630];
    end
    always @(spike_out_source_array[631]) begin 
        spike_out_source631 = spike_out_source_array[631];
    end
    always @(spike_out_source_array[632]) begin 
        spike_out_source632 = spike_out_source_array[632];
    end
    always @(spike_out_source_array[633]) begin 
        spike_out_source633 = spike_out_source_array[633];
    end
    always @(spike_out_source_array[634]) begin 
        spike_out_source634 = spike_out_source_array[634];
    end
    always @(spike_out_source_array[635]) begin 
        spike_out_source635 = spike_out_source_array[635];
    end
    always @(spike_out_source_array[636]) begin 
        spike_out_source636 = spike_out_source_array[636];
    end
    always @(spike_out_source_array[637]) begin 
        spike_out_source637 = spike_out_source_array[637];
    end
    always @(spike_out_source_array[638]) begin 
        spike_out_source638 = spike_out_source_array[638];
    end
    always @(spike_out_source_array[639]) begin 
        spike_out_source639 = spike_out_source_array[639];
    end
    always @(spike_out_source_array[640]) begin 
        spike_out_source640 = spike_out_source_array[640];
    end
    always @(spike_out_source_array[641]) begin 
        spike_out_source641 = spike_out_source_array[641];
    end
    always @(spike_out_source_array[642]) begin 
        spike_out_source642 = spike_out_source_array[642];
    end
    always @(spike_out_source_array[643]) begin 
        spike_out_source643 = spike_out_source_array[643];
    end
    always @(spike_out_source_array[644]) begin 
        spike_out_source644 = spike_out_source_array[644];
    end
    always @(spike_out_source_array[645]) begin 
        spike_out_source645 = spike_out_source_array[645];
    end
    always @(spike_out_source_array[646]) begin 
        spike_out_source646 = spike_out_source_array[646];
    end
    always @(spike_out_source_array[647]) begin 
        spike_out_source647 = spike_out_source_array[647];
    end
    always @(spike_out_source_array[648]) begin 
        spike_out_source648 = spike_out_source_array[648];
    end
    always @(spike_out_source_array[649]) begin 
        spike_out_source649 = spike_out_source_array[649];
    end
    always @(spike_out_source_array[650]) begin 
        spike_out_source650 = spike_out_source_array[650];
    end
    always @(spike_out_source_array[651]) begin 
        spike_out_source651 = spike_out_source_array[651];
    end
    always @(spike_out_source_array[652]) begin 
        spike_out_source652 = spike_out_source_array[652];
    end
    always @(spike_out_source_array[653]) begin 
        spike_out_source653 = spike_out_source_array[653];
    end
    always @(spike_out_source_array[654]) begin 
        spike_out_source654 = spike_out_source_array[654];
    end
    always @(spike_out_source_array[655]) begin 
        spike_out_source655 = spike_out_source_array[655];
    end
    always @(spike_out_source_array[656]) begin 
        spike_out_source656 = spike_out_source_array[656];
    end
    always @(spike_out_source_array[657]) begin 
        spike_out_source657 = spike_out_source_array[657];
    end
    always @(spike_out_source_array[658]) begin 
        spike_out_source658 = spike_out_source_array[658];
    end
    always @(spike_out_source_array[659]) begin 
        spike_out_source659 = spike_out_source_array[659];
    end
    always @(spike_out_source_array[660]) begin 
        spike_out_source660 = spike_out_source_array[660];
    end
    always @(spike_out_source_array[661]) begin 
        spike_out_source661 = spike_out_source_array[661];
    end
    always @(spike_out_source_array[662]) begin 
        spike_out_source662 = spike_out_source_array[662];
    end
    always @(spike_out_source_array[663]) begin 
        spike_out_source663 = spike_out_source_array[663];
    end
    always @(spike_out_source_array[664]) begin 
        spike_out_source664 = spike_out_source_array[664];
    end
    always @(spike_out_source_array[665]) begin 
        spike_out_source665 = spike_out_source_array[665];
    end
    always @(spike_out_source_array[666]) begin 
        spike_out_source666 = spike_out_source_array[666];
    end
    always @(spike_out_source_array[667]) begin 
        spike_out_source667 = spike_out_source_array[667];
    end
    always @(spike_out_source_array[668]) begin 
        spike_out_source668 = spike_out_source_array[668];
    end
    always @(spike_out_source_array[669]) begin 
        spike_out_source669 = spike_out_source_array[669];
    end
    always @(spike_out_source_array[670]) begin 
        spike_out_source670 = spike_out_source_array[670];
    end
    always @(spike_out_source_array[671]) begin 
        spike_out_source671 = spike_out_source_array[671];
    end
    always @(spike_out_source_array[672]) begin 
        spike_out_source672 = spike_out_source_array[672];
    end
    always @(spike_out_source_array[673]) begin 
        spike_out_source673 = spike_out_source_array[673];
    end
    always @(spike_out_source_array[674]) begin 
        spike_out_source674 = spike_out_source_array[674];
    end
    always @(spike_out_source_array[675]) begin 
        spike_out_source675 = spike_out_source_array[675];
    end
    always @(spike_out_source_array[676]) begin 
        spike_out_source676 = spike_out_source_array[676];
    end
    always @(spike_out_source_array[677]) begin 
        spike_out_source677 = spike_out_source_array[677];
    end
    always @(spike_out_source_array[678]) begin 
        spike_out_source678 = spike_out_source_array[678];
    end
    always @(spike_out_source_array[679]) begin 
        spike_out_source679 = spike_out_source_array[679];
    end
    always @(spike_out_source_array[680]) begin 
        spike_out_source680 = spike_out_source_array[680];
    end
    always @(spike_out_source_array[681]) begin 
        spike_out_source681 = spike_out_source_array[681];
    end
    always @(spike_out_source_array[682]) begin 
        spike_out_source682 = spike_out_source_array[682];
    end
    always @(spike_out_source_array[683]) begin 
        spike_out_source683 = spike_out_source_array[683];
    end
    always @(spike_out_source_array[684]) begin 
        spike_out_source684 = spike_out_source_array[684];
    end
    always @(spike_out_source_array[685]) begin 
        spike_out_source685 = spike_out_source_array[685];
    end
    always @(spike_out_source_array[686]) begin 
        spike_out_source686 = spike_out_source_array[686];
    end
    always @(spike_out_source_array[687]) begin 
        spike_out_source687 = spike_out_source_array[687];
    end
    always @(spike_out_source_array[688]) begin 
        spike_out_source688 = spike_out_source_array[688];
    end
    always @(spike_out_source_array[689]) begin 
        spike_out_source689 = spike_out_source_array[689];
    end
    always @(spike_out_source_array[690]) begin 
        spike_out_source690 = spike_out_source_array[690];
    end
    always @(spike_out_source_array[691]) begin 
        spike_out_source691 = spike_out_source_array[691];
    end
    always @(spike_out_source_array[692]) begin 
        spike_out_source692 = spike_out_source_array[692];
    end
    always @(spike_out_source_array[693]) begin 
        spike_out_source693 = spike_out_source_array[693];
    end
    always @(spike_out_source_array[694]) begin 
        spike_out_source694 = spike_out_source_array[694];
    end
    always @(spike_out_source_array[695]) begin 
        spike_out_source695 = spike_out_source_array[695];
    end
    always @(spike_out_source_array[696]) begin 
        spike_out_source696 = spike_out_source_array[696];
    end
    always @(spike_out_source_array[697]) begin 
        spike_out_source697 = spike_out_source_array[697];
    end
    always @(spike_out_source_array[698]) begin 
        spike_out_source698 = spike_out_source_array[698];
    end
    always @(spike_out_source_array[699]) begin 
        spike_out_source699 = spike_out_source_array[699];
    end
    always @(spike_out_source_array[700]) begin 
        spike_out_source700 = spike_out_source_array[700];
    end
    always @(spike_out_source_array[701]) begin 
        spike_out_source701 = spike_out_source_array[701];
    end
    always @(spike_out_source_array[702]) begin 
        spike_out_source702 = spike_out_source_array[702];
    end
    always @(spike_out_source_array[703]) begin 
        spike_out_source703 = spike_out_source_array[703];
    end
    always @(spike_out_source_array[704]) begin 
        spike_out_source704 = spike_out_source_array[704];
    end
    always @(spike_out_source_array[705]) begin 
        spike_out_source705 = spike_out_source_array[705];
    end
    always @(spike_out_source_array[706]) begin 
        spike_out_source706 = spike_out_source_array[706];
    end
    always @(spike_out_source_array[707]) begin 
        spike_out_source707 = spike_out_source_array[707];
    end
    always @(spike_out_source_array[708]) begin 
        spike_out_source708 = spike_out_source_array[708];
    end
    always @(spike_out_source_array[709]) begin 
        spike_out_source709 = spike_out_source_array[709];
    end
    always @(spike_out_source_array[710]) begin 
        spike_out_source710 = spike_out_source_array[710];
    end
    always @(spike_out_source_array[711]) begin 
        spike_out_source711 = spike_out_source_array[711];
    end
    always @(spike_out_source_array[712]) begin 
        spike_out_source712 = spike_out_source_array[712];
    end
    always @(spike_out_source_array[713]) begin 
        spike_out_source713 = spike_out_source_array[713];
    end
    always @(spike_out_source_array[714]) begin 
        spike_out_source714 = spike_out_source_array[714];
    end
    always @(spike_out_source_array[715]) begin 
        spike_out_source715 = spike_out_source_array[715];
    end
    always @(spike_out_source_array[716]) begin 
        spike_out_source716 = spike_out_source_array[716];
    end
    always @(spike_out_source_array[717]) begin 
        spike_out_source717 = spike_out_source_array[717];
    end
    always @(spike_out_source_array[718]) begin 
        spike_out_source718 = spike_out_source_array[718];
    end
    always @(spike_out_source_array[719]) begin 
        spike_out_source719 = spike_out_source_array[719];
    end
    always @(spike_out_source_array[720]) begin 
        spike_out_source720 = spike_out_source_array[720];
    end
    always @(spike_out_source_array[721]) begin 
        spike_out_source721 = spike_out_source_array[721];
    end
    always @(spike_out_source_array[722]) begin 
        spike_out_source722 = spike_out_source_array[722];
    end
    always @(spike_out_source_array[723]) begin 
        spike_out_source723 = spike_out_source_array[723];
    end
    always @(spike_out_source_array[724]) begin 
        spike_out_source724 = spike_out_source_array[724];
    end
    always @(spike_out_source_array[725]) begin 
        spike_out_source725 = spike_out_source_array[725];
    end
    always @(spike_out_source_array[726]) begin 
        spike_out_source726 = spike_out_source_array[726];
    end
    always @(spike_out_source_array[727]) begin 
        spike_out_source727 = spike_out_source_array[727];
    end
    always @(spike_out_source_array[728]) begin 
        spike_out_source728 = spike_out_source_array[728];
    end
    always @(spike_out_source_array[729]) begin 
        spike_out_source729 = spike_out_source_array[729];
    end
    always @(spike_out_source_array[730]) begin 
        spike_out_source730 = spike_out_source_array[730];
    end
    always @(spike_out_source_array[731]) begin 
        spike_out_source731 = spike_out_source_array[731];
    end
    always @(spike_out_source_array[732]) begin 
        spike_out_source732 = spike_out_source_array[732];
    end
    always @(spike_out_source_array[733]) begin 
        spike_out_source733 = spike_out_source_array[733];
    end
    always @(spike_out_source_array[734]) begin 
        spike_out_source734 = spike_out_source_array[734];
    end
    always @(spike_out_source_array[735]) begin 
        spike_out_source735 = spike_out_source_array[735];
    end
    always @(spike_out_source_array[736]) begin 
        spike_out_source736 = spike_out_source_array[736];
    end
    always @(spike_out_source_array[737]) begin 
        spike_out_source737 = spike_out_source_array[737];
    end
    always @(spike_out_source_array[738]) begin 
        spike_out_source738 = spike_out_source_array[738];
    end
    always @(spike_out_source_array[739]) begin 
        spike_out_source739 = spike_out_source_array[739];
    end
    always @(spike_out_source_array[740]) begin 
        spike_out_source740 = spike_out_source_array[740];
    end
    always @(spike_out_source_array[741]) begin 
        spike_out_source741 = spike_out_source_array[741];
    end
    always @(spike_out_source_array[742]) begin 
        spike_out_source742 = spike_out_source_array[742];
    end
    always @(spike_out_source_array[743]) begin 
        spike_out_source743 = spike_out_source_array[743];
    end
    always @(spike_out_source_array[744]) begin 
        spike_out_source744 = spike_out_source_array[744];
    end
    always @(spike_out_source_array[745]) begin 
        spike_out_source745 = spike_out_source_array[745];
    end
    always @(spike_out_source_array[746]) begin 
        spike_out_source746 = spike_out_source_array[746];
    end
    always @(spike_out_source_array[747]) begin 
        spike_out_source747 = spike_out_source_array[747];
    end
    always @(spike_out_source_array[748]) begin 
        spike_out_source748 = spike_out_source_array[748];
    end
    always @(spike_out_source_array[749]) begin 
        spike_out_source749 = spike_out_source_array[749];
    end
    always @(spike_out_source_array[750]) begin 
        spike_out_source750 = spike_out_source_array[750];
    end
    always @(spike_out_source_array[751]) begin 
        spike_out_source751 = spike_out_source_array[751];
    end
    always @(spike_out_source_array[752]) begin 
        spike_out_source752 = spike_out_source_array[752];
    end
    always @(spike_out_source_array[753]) begin 
        spike_out_source753 = spike_out_source_array[753];
    end
    always @(spike_out_source_array[754]) begin 
        spike_out_source754 = spike_out_source_array[754];
    end
    always @(spike_out_source_array[755]) begin 
        spike_out_source755 = spike_out_source_array[755];
    end
    always @(spike_out_source_array[756]) begin 
        spike_out_source756 = spike_out_source_array[756];
    end
    always @(spike_out_source_array[757]) begin 
        spike_out_source757 = spike_out_source_array[757];
    end
    always @(spike_out_source_array[758]) begin 
        spike_out_source758 = spike_out_source_array[758];
    end
    always @(spike_out_source_array[759]) begin 
        spike_out_source759 = spike_out_source_array[759];
    end
    always @(spike_out_source_array[760]) begin 
        spike_out_source760 = spike_out_source_array[760];
    end
    always @(spike_out_source_array[761]) begin 
        spike_out_source761 = spike_out_source_array[761];
    end
    always @(spike_out_source_array[762]) begin 
        spike_out_source762 = spike_out_source_array[762];
    end
    always @(spike_out_source_array[763]) begin 
        spike_out_source763 = spike_out_source_array[763];
    end
    always @(spike_out_source_array[764]) begin 
        spike_out_source764 = spike_out_source_array[764];
    end
    always @(spike_out_source_array[765]) begin 
        spike_out_source765 = spike_out_source_array[765];
    end
    always @(spike_out_source_array[766]) begin 
        spike_out_source766 = spike_out_source_array[766];
    end
    always @(spike_out_source_array[767]) begin 
        spike_out_source767 = spike_out_source_array[767];
    end
    always @(spike_out_source_array[768]) begin 
        spike_out_source768 = spike_out_source_array[768];
    end
    always @(spike_out_source_array[769]) begin 
        spike_out_source769 = spike_out_source_array[769];
    end
    always @(spike_out_source_array[770]) begin 
        spike_out_source770 = spike_out_source_array[770];
    end
    always @(spike_out_source_array[771]) begin 
        spike_out_source771 = spike_out_source_array[771];
    end
    always @(spike_out_source_array[772]) begin 
        spike_out_source772 = spike_out_source_array[772];
    end
    always @(spike_out_source_array[773]) begin 
        spike_out_source773 = spike_out_source_array[773];
    end
    always @(spike_out_source_array[774]) begin 
        spike_out_source774 = spike_out_source_array[774];
    end
    always @(spike_out_source_array[775]) begin 
        spike_out_source775 = spike_out_source_array[775];
    end
    always @(spike_out_source_array[776]) begin 
        spike_out_source776 = spike_out_source_array[776];
    end
    always @(spike_out_source_array[777]) begin 
        spike_out_source777 = spike_out_source_array[777];
    end
    always @(spike_out_source_array[778]) begin 
        spike_out_source778 = spike_out_source_array[778];
    end
    always @(spike_out_source_array[779]) begin 
        spike_out_source779 = spike_out_source_array[779];
    end
    always @(spike_out_source_array[780]) begin 
        spike_out_source780 = spike_out_source_array[780];
    end
    always @(spike_out_source_array[781]) begin 
        spike_out_source781 = spike_out_source_array[781];
    end
    always @(spike_out_source_array[782]) begin 
        spike_out_source782 = spike_out_source_array[782];
    end
    always @(spike_out_source_array[783]) begin 
        spike_out_source783 = spike_out_source_array[783];
    end
    always @(spike_out_source_array[784]) begin 
        spike_out_source784 = spike_out_source_array[784];
    end
    always @(spike_out_source_array[785]) begin 
        spike_out_source785 = spike_out_source_array[785];
    end
    always @(spike_out_source_array[786]) begin 
        spike_out_source786 = spike_out_source_array[786];
    end
    always @(spike_out_source_array[787]) begin 
        spike_out_source787 = spike_out_source_array[787];
    end
    always @(spike_out_source_array[788]) begin 
        spike_out_source788 = spike_out_source_array[788];
    end
    always @(spike_out_source_array[789]) begin 
        spike_out_source789 = spike_out_source_array[789];
    end
    always @(spike_out_source_array[790]) begin 
        spike_out_source790 = spike_out_source_array[790];
    end
    always @(spike_out_source_array[791]) begin 
        spike_out_source791 = spike_out_source_array[791];
    end
    always @(spike_out_source_array[792]) begin 
        spike_out_source792 = spike_out_source_array[792];
    end
    always @(spike_out_source_array[793]) begin 
        spike_out_source793 = spike_out_source_array[793];
    end
    always @(spike_out_source_array[794]) begin 
        spike_out_source794 = spike_out_source_array[794];
    end
    always @(spike_out_source_array[795]) begin 
        spike_out_source795 = spike_out_source_array[795];
    end
    always @(spike_out_source_array[796]) begin 
        spike_out_source796 = spike_out_source_array[796];
    end
    always @(spike_out_source_array[797]) begin 
        spike_out_source797 = spike_out_source_array[797];
    end
    always @(spike_out_source_array[798]) begin 
        spike_out_source798 = spike_out_source_array[798];
    end
    always @(spike_out_source_array[799]) begin 
        spike_out_source799 = spike_out_source_array[799];
    end
    always @(spike_out_source_array[800]) begin 
        spike_out_source800 = spike_out_source_array[800];
    end
    always @(spike_out_source_array[801]) begin 
        spike_out_source801 = spike_out_source_array[801];
    end
    always @(spike_out_source_array[802]) begin 
        spike_out_source802 = spike_out_source_array[802];
    end
    always @(spike_out_source_array[803]) begin 
        spike_out_source803 = spike_out_source_array[803];
    end
    always @(spike_out_source_array[804]) begin 
        spike_out_source804 = spike_out_source_array[804];
    end
    always @(spike_out_source_array[805]) begin 
        spike_out_source805 = spike_out_source_array[805];
    end
    always @(spike_out_source_array[806]) begin 
        spike_out_source806 = spike_out_source_array[806];
    end
    always @(spike_out_source_array[807]) begin 
        spike_out_source807 = spike_out_source_array[807];
    end
    always @(spike_out_source_array[808]) begin 
        spike_out_source808 = spike_out_source_array[808];
    end
    always @(spike_out_source_array[809]) begin 
        spike_out_source809 = spike_out_source_array[809];
    end
    always @(spike_out_source_array[810]) begin 
        spike_out_source810 = spike_out_source_array[810];
    end
    always @(spike_out_source_array[811]) begin 
        spike_out_source811 = spike_out_source_array[811];
    end
    always @(spike_out_source_array[812]) begin 
        spike_out_source812 = spike_out_source_array[812];
    end
    always @(spike_out_source_array[813]) begin 
        spike_out_source813 = spike_out_source_array[813];
    end
    always @(spike_out_source_array[814]) begin 
        spike_out_source814 = spike_out_source_array[814];
    end
    always @(spike_out_source_array[815]) begin 
        spike_out_source815 = spike_out_source_array[815];
    end
    always @(spike_out_source_array[816]) begin 
        spike_out_source816 = spike_out_source_array[816];
    end
    always @(spike_out_source_array[817]) begin 
        spike_out_source817 = spike_out_source_array[817];
    end
    always @(spike_out_source_array[818]) begin 
        spike_out_source818 = spike_out_source_array[818];
    end
    always @(spike_out_source_array[819]) begin 
        spike_out_source819 = spike_out_source_array[819];
    end
    always @(spike_out_source_array[820]) begin 
        spike_out_source820 = spike_out_source_array[820];
    end
    always @(spike_out_source_array[821]) begin 
        spike_out_source821 = spike_out_source_array[821];
    end
    always @(spike_out_source_array[822]) begin 
        spike_out_source822 = spike_out_source_array[822];
    end
    always @(spike_out_source_array[823]) begin 
        spike_out_source823 = spike_out_source_array[823];
    end
    always @(spike_out_source_array[824]) begin 
        spike_out_source824 = spike_out_source_array[824];
    end
    always @(spike_out_source_array[825]) begin 
        spike_out_source825 = spike_out_source_array[825];
    end
    always @(spike_out_source_array[826]) begin 
        spike_out_source826 = spike_out_source_array[826];
    end
    always @(spike_out_source_array[827]) begin 
        spike_out_source827 = spike_out_source_array[827];
    end
    always @(spike_out_source_array[828]) begin 
        spike_out_source828 = spike_out_source_array[828];
    end
    always @(spike_out_source_array[829]) begin 
        spike_out_source829 = spike_out_source_array[829];
    end
    always @(spike_out_source_array[830]) begin 
        spike_out_source830 = spike_out_source_array[830];
    end
    always @(spike_out_source_array[831]) begin 
        spike_out_source831 = spike_out_source_array[831];
    end
    always @(spike_out_source_array[832]) begin 
        spike_out_source832 = spike_out_source_array[832];
    end
    always @(spike_out_source_array[833]) begin 
        spike_out_source833 = spike_out_source_array[833];
    end
    always @(spike_out_source_array[834]) begin 
        spike_out_source834 = spike_out_source_array[834];
    end
    always @(spike_out_source_array[835]) begin 
        spike_out_source835 = spike_out_source_array[835];
    end
    always @(spike_out_source_array[836]) begin 
        spike_out_source836 = spike_out_source_array[836];
    end
    always @(spike_out_source_array[837]) begin 
        spike_out_source837 = spike_out_source_array[837];
    end
    always @(spike_out_source_array[838]) begin 
        spike_out_source838 = spike_out_source_array[838];
    end
    always @(spike_out_source_array[839]) begin 
        spike_out_source839 = spike_out_source_array[839];
    end
    always @(spike_out_source_array[840]) begin 
        spike_out_source840 = spike_out_source_array[840];
    end
    always @(spike_out_source_array[841]) begin 
        spike_out_source841 = spike_out_source_array[841];
    end
    always @(spike_out_source_array[842]) begin 
        spike_out_source842 = spike_out_source_array[842];
    end
    always @(spike_out_source_array[843]) begin 
        spike_out_source843 = spike_out_source_array[843];
    end
    always @(spike_out_source_array[844]) begin 
        spike_out_source844 = spike_out_source_array[844];
    end
    always @(spike_out_source_array[845]) begin 
        spike_out_source845 = spike_out_source_array[845];
    end
    always @(spike_out_source_array[846]) begin 
        spike_out_source846 = spike_out_source_array[846];
    end
    always @(spike_out_source_array[847]) begin 
        spike_out_source847 = spike_out_source_array[847];
    end
    always @(spike_out_source_array[848]) begin 
        spike_out_source848 = spike_out_source_array[848];
    end
    always @(spike_out_source_array[849]) begin 
        spike_out_source849 = spike_out_source_array[849];
    end
    always @(spike_out_source_array[850]) begin 
        spike_out_source850 = spike_out_source_array[850];
    end
    always @(spike_out_source_array[851]) begin 
        spike_out_source851 = spike_out_source_array[851];
    end
    always @(spike_out_source_array[852]) begin 
        spike_out_source852 = spike_out_source_array[852];
    end
    always @(spike_out_source_array[853]) begin 
        spike_out_source853 = spike_out_source_array[853];
    end
    always @(spike_out_source_array[854]) begin 
        spike_out_source854 = spike_out_source_array[854];
    end
    always @(spike_out_source_array[855]) begin 
        spike_out_source855 = spike_out_source_array[855];
    end
    always @(spike_out_source_array[856]) begin 
        spike_out_source856 = spike_out_source_array[856];
    end
    always @(spike_out_source_array[857]) begin 
        spike_out_source857 = spike_out_source_array[857];
    end
    always @(spike_out_source_array[858]) begin 
        spike_out_source858 = spike_out_source_array[858];
    end
    always @(spike_out_source_array[859]) begin 
        spike_out_source859 = spike_out_source_array[859];
    end
    always @(spike_out_source_array[860]) begin 
        spike_out_source860 = spike_out_source_array[860];
    end
    always @(spike_out_source_array[861]) begin 
        spike_out_source861 = spike_out_source_array[861];
    end
    always @(spike_out_source_array[862]) begin 
        spike_out_source862 = spike_out_source_array[862];
    end
    always @(spike_out_source_array[863]) begin 
        spike_out_source863 = spike_out_source_array[863];
    end
    always @(spike_out_source_array[864]) begin 
        spike_out_source864 = spike_out_source_array[864];
    end
    always @(spike_out_source_array[865]) begin 
        spike_out_source865 = spike_out_source_array[865];
    end
    always @(spike_out_source_array[866]) begin 
        spike_out_source866 = spike_out_source_array[866];
    end
    always @(spike_out_source_array[867]) begin 
        spike_out_source867 = spike_out_source_array[867];
    end
    always @(spike_out_source_array[868]) begin 
        spike_out_source868 = spike_out_source_array[868];
    end
    always @(spike_out_source_array[869]) begin 
        spike_out_source869 = spike_out_source_array[869];
    end
    always @(spike_out_source_array[870]) begin 
        spike_out_source870 = spike_out_source_array[870];
    end
    always @(spike_out_source_array[871]) begin 
        spike_out_source871 = spike_out_source_array[871];
    end
    always @(spike_out_source_array[872]) begin 
        spike_out_source872 = spike_out_source_array[872];
    end
    always @(spike_out_source_array[873]) begin 
        spike_out_source873 = spike_out_source_array[873];
    end
    always @(spike_out_source_array[874]) begin 
        spike_out_source874 = spike_out_source_array[874];
    end
    always @(spike_out_source_array[875]) begin 
        spike_out_source875 = spike_out_source_array[875];
    end
    always @(spike_out_source_array[876]) begin 
        spike_out_source876 = spike_out_source_array[876];
    end
    always @(spike_out_source_array[877]) begin 
        spike_out_source877 = spike_out_source_array[877];
    end
    always @(spike_out_source_array[878]) begin 
        spike_out_source878 = spike_out_source_array[878];
    end
    always @(spike_out_source_array[879]) begin 
        spike_out_source879 = spike_out_source_array[879];
    end
    always @(spike_out_source_array[880]) begin 
        spike_out_source880 = spike_out_source_array[880];
    end
    always @(spike_out_source_array[881]) begin 
        spike_out_source881 = spike_out_source_array[881];
    end
    always @(spike_out_source_array[882]) begin 
        spike_out_source882 = spike_out_source_array[882];
    end
    always @(spike_out_source_array[883]) begin 
        spike_out_source883 = spike_out_source_array[883];
    end
    always @(spike_out_source_array[884]) begin 
        spike_out_source884 = spike_out_source_array[884];
    end
    always @(spike_out_source_array[885]) begin 
        spike_out_source885 = spike_out_source_array[885];
    end
    always @(spike_out_source_array[886]) begin 
        spike_out_source886 = spike_out_source_array[886];
    end
    always @(spike_out_source_array[887]) begin 
        spike_out_source887 = spike_out_source_array[887];
    end
    always @(spike_out_source_array[888]) begin 
        spike_out_source888 = spike_out_source_array[888];
    end
    always @(spike_out_source_array[889]) begin 
        spike_out_source889 = spike_out_source_array[889];
    end
    always @(spike_out_source_array[890]) begin 
        spike_out_source890 = spike_out_source_array[890];
    end
    always @(spike_out_source_array[891]) begin 
        spike_out_source891 = spike_out_source_array[891];
    end
    always @(spike_out_source_array[892]) begin 
        spike_out_source892 = spike_out_source_array[892];
    end
    always @(spike_out_source_array[893]) begin 
        spike_out_source893 = spike_out_source_array[893];
    end
    always @(spike_out_source_array[894]) begin 
        spike_out_source894 = spike_out_source_array[894];
    end
    always @(spike_out_source_array[895]) begin 
        spike_out_source895 = spike_out_source_array[895];
    end
    always @(spike_out_source_array[896]) begin 
        spike_out_source896 = spike_out_source_array[896];
    end
    always @(spike_out_source_array[897]) begin 
        spike_out_source897 = spike_out_source_array[897];
    end
    always @(spike_out_source_array[898]) begin 
        spike_out_source898 = spike_out_source_array[898];
    end
    always @(spike_out_source_array[899]) begin 
        spike_out_source899 = spike_out_source_array[899];
    end
    always @(spike_out_source_array[900]) begin 
        spike_out_source900 = spike_out_source_array[900];
    end
    always @(spike_out_source_array[901]) begin 
        spike_out_source901 = spike_out_source_array[901];
    end
    always @(spike_out_source_array[902]) begin 
        spike_out_source902 = spike_out_source_array[902];
    end
    always @(spike_out_source_array[903]) begin 
        spike_out_source903 = spike_out_source_array[903];
    end
    always @(spike_out_source_array[904]) begin 
        spike_out_source904 = spike_out_source_array[904];
    end
    always @(spike_out_source_array[905]) begin 
        spike_out_source905 = spike_out_source_array[905];
    end
    always @(spike_out_source_array[906]) begin 
        spike_out_source906 = spike_out_source_array[906];
    end
    always @(spike_out_source_array[907]) begin 
        spike_out_source907 = spike_out_source_array[907];
    end
    always @(spike_out_source_array[908]) begin 
        spike_out_source908 = spike_out_source_array[908];
    end
    always @(spike_out_source_array[909]) begin 
        spike_out_source909 = spike_out_source_array[909];
    end
    always @(spike_out_source_array[910]) begin 
        spike_out_source910 = spike_out_source_array[910];
    end
    always @(spike_out_source_array[911]) begin 
        spike_out_source911 = spike_out_source_array[911];
    end
    always @(spike_out_source_array[912]) begin 
        spike_out_source912 = spike_out_source_array[912];
    end
    always @(spike_out_source_array[913]) begin 
        spike_out_source913 = spike_out_source_array[913];
    end
    always @(spike_out_source_array[914]) begin 
        spike_out_source914 = spike_out_source_array[914];
    end
    always @(spike_out_source_array[915]) begin 
        spike_out_source915 = spike_out_source_array[915];
    end
    always @(spike_out_source_array[916]) begin 
        spike_out_source916 = spike_out_source_array[916];
    end
    always @(spike_out_source_array[917]) begin 
        spike_out_source917 = spike_out_source_array[917];
    end
    always @(spike_out_source_array[918]) begin 
        spike_out_source918 = spike_out_source_array[918];
    end
    always @(spike_out_source_array[919]) begin 
        spike_out_source919 = spike_out_source_array[919];
    end
    always @(spike_out_source_array[920]) begin 
        spike_out_source920 = spike_out_source_array[920];
    end
    always @(spike_out_source_array[921]) begin 
        spike_out_source921 = spike_out_source_array[921];
    end
    always @(spike_out_source_array[922]) begin 
        spike_out_source922 = spike_out_source_array[922];
    end
    always @(spike_out_source_array[923]) begin 
        spike_out_source923 = spike_out_source_array[923];
    end
    always @(spike_out_source_array[924]) begin 
        spike_out_source924 = spike_out_source_array[924];
    end
    always @(spike_out_source_array[925]) begin 
        spike_out_source925 = spike_out_source_array[925];
    end
    always @(spike_out_source_array[926]) begin 
        spike_out_source926 = spike_out_source_array[926];
    end
    always @(spike_out_source_array[927]) begin 
        spike_out_source927 = spike_out_source_array[927];
    end
    always @(spike_out_source_array[928]) begin 
        spike_out_source928 = spike_out_source_array[928];
    end
    always @(spike_out_source_array[929]) begin 
        spike_out_source929 = spike_out_source_array[929];
    end
    always @(spike_out_source_array[930]) begin 
        spike_out_source930 = spike_out_source_array[930];
    end
    always @(spike_out_source_array[931]) begin 
        spike_out_source931 = spike_out_source_array[931];
    end
    always @(spike_out_source_array[932]) begin 
        spike_out_source932 = spike_out_source_array[932];
    end
    always @(spike_out_source_array[933]) begin 
        spike_out_source933 = spike_out_source_array[933];
    end
    always @(spike_out_source_array[934]) begin 
        spike_out_source934 = spike_out_source_array[934];
    end
    always @(spike_out_source_array[935]) begin 
        spike_out_source935 = spike_out_source_array[935];
    end
    always @(spike_out_source_array[936]) begin 
        spike_out_source936 = spike_out_source_array[936];
    end
    always @(spike_out_source_array[937]) begin 
        spike_out_source937 = spike_out_source_array[937];
    end
    always @(spike_out_source_array[938]) begin 
        spike_out_source938 = spike_out_source_array[938];
    end
    always @(spike_out_source_array[939]) begin 
        spike_out_source939 = spike_out_source_array[939];
    end
    always @(spike_out_source_array[940]) begin 
        spike_out_source940 = spike_out_source_array[940];
    end
    always @(spike_out_source_array[941]) begin 
        spike_out_source941 = spike_out_source_array[941];
    end
    always @(spike_out_source_array[942]) begin 
        spike_out_source942 = spike_out_source_array[942];
    end
    always @(spike_out_source_array[943]) begin 
        spike_out_source943 = spike_out_source_array[943];
    end
    always @(spike_out_source_array[944]) begin 
        spike_out_source944 = spike_out_source_array[944];
    end
    always @(spike_out_source_array[945]) begin 
        spike_out_source945 = spike_out_source_array[945];
    end
    always @(spike_out_source_array[946]) begin 
        spike_out_source946 = spike_out_source_array[946];
    end
    always @(spike_out_source_array[947]) begin 
        spike_out_source947 = spike_out_source_array[947];
    end
    always @(spike_out_source_array[948]) begin 
        spike_out_source948 = spike_out_source_array[948];
    end
    always @(spike_out_source_array[949]) begin 
        spike_out_source949 = spike_out_source_array[949];
    end
    always @(spike_out_source_array[950]) begin 
        spike_out_source950 = spike_out_source_array[950];
    end
    always @(spike_out_source_array[951]) begin 
        spike_out_source951 = spike_out_source_array[951];
    end
    always @(spike_out_source_array[952]) begin 
        spike_out_source952 = spike_out_source_array[952];
    end
    always @(spike_out_source_array[953]) begin 
        spike_out_source953 = spike_out_source_array[953];
    end
    always @(spike_out_source_array[954]) begin 
        spike_out_source954 = spike_out_source_array[954];
    end
    always @(spike_out_source_array[955]) begin 
        spike_out_source955 = spike_out_source_array[955];
    end
    always @(spike_out_source_array[956]) begin 
        spike_out_source956 = spike_out_source_array[956];
    end
    always @(spike_out_source_array[957]) begin 
        spike_out_source957 = spike_out_source_array[957];
    end
    always @(spike_out_source_array[958]) begin 
        spike_out_source958 = spike_out_source_array[958];
    end
    always @(spike_out_source_array[959]) begin 
        spike_out_source959 = spike_out_source_array[959];
    end
    always @(spike_out_source_array[960]) begin 
        spike_out_source960 = spike_out_source_array[960];
    end
    always @(spike_out_source_array[961]) begin 
        spike_out_source961 = spike_out_source_array[961];
    end
    always @(spike_out_source_array[962]) begin 
        spike_out_source962 = spike_out_source_array[962];
    end
    always @(spike_out_source_array[963]) begin 
        spike_out_source963 = spike_out_source_array[963];
    end
    always @(spike_out_source_array[964]) begin 
        spike_out_source964 = spike_out_source_array[964];
    end
    always @(spike_out_source_array[965]) begin 
        spike_out_source965 = spike_out_source_array[965];
    end
    always @(spike_out_source_array[966]) begin 
        spike_out_source966 = spike_out_source_array[966];
    end
    always @(spike_out_source_array[967]) begin 
        spike_out_source967 = spike_out_source_array[967];
    end
    always @(spike_out_source_array[968]) begin 
        spike_out_source968 = spike_out_source_array[968];
    end
    always @(spike_out_source_array[969]) begin 
        spike_out_source969 = spike_out_source_array[969];
    end
    always @(spike_out_source_array[970]) begin 
        spike_out_source970 = spike_out_source_array[970];
    end
    always @(spike_out_source_array[971]) begin 
        spike_out_source971 = spike_out_source_array[971];
    end
    always @(spike_out_source_array[972]) begin 
        spike_out_source972 = spike_out_source_array[972];
    end
    always @(spike_out_source_array[973]) begin 
        spike_out_source973 = spike_out_source_array[973];
    end
    always @(spike_out_source_array[974]) begin 
        spike_out_source974 = spike_out_source_array[974];
    end
    always @(spike_out_source_array[975]) begin 
        spike_out_source975 = spike_out_source_array[975];
    end
    always @(spike_out_source_array[976]) begin 
        spike_out_source976 = spike_out_source_array[976];
    end
    always @(spike_out_source_array[977]) begin 
        spike_out_source977 = spike_out_source_array[977];
    end
    always @(spike_out_source_array[978]) begin 
        spike_out_source978 = spike_out_source_array[978];
    end
    always @(spike_out_source_array[979]) begin 
        spike_out_source979 = spike_out_source_array[979];
    end
    always @(spike_out_source_array[980]) begin 
        spike_out_source980 = spike_out_source_array[980];
    end
    always @(spike_out_source_array[981]) begin 
        spike_out_source981 = spike_out_source_array[981];
    end
    always @(spike_out_source_array[982]) begin 
        spike_out_source982 = spike_out_source_array[982];
    end
    always @(spike_out_source_array[983]) begin 
        spike_out_source983 = spike_out_source_array[983];
    end
    always @(spike_out_source_array[984]) begin 
        spike_out_source984 = spike_out_source_array[984];
    end
    always @(spike_out_source_array[985]) begin 
        spike_out_source985 = spike_out_source_array[985];
    end
    always @(spike_out_source_array[986]) begin 
        spike_out_source986 = spike_out_source_array[986];
    end
    always @(spike_out_source_array[987]) begin 
        spike_out_source987 = spike_out_source_array[987];
    end
    always @(spike_out_source_array[988]) begin 
        spike_out_source988 = spike_out_source_array[988];
    end
    always @(spike_out_source_array[989]) begin 
        spike_out_source989 = spike_out_source_array[989];
    end
    always @(spike_out_source_array[990]) begin 
        spike_out_source990 = spike_out_source_array[990];
    end
    always @(spike_out_source_array[991]) begin 
        spike_out_source991 = spike_out_source_array[991];
    end
    always @(spike_out_source_array[992]) begin 
        spike_out_source992 = spike_out_source_array[992];
    end
    always @(spike_out_source_array[993]) begin 
        spike_out_source993 = spike_out_source_array[993];
    end
    always @(spike_out_source_array[994]) begin 
        spike_out_source994 = spike_out_source_array[994];
    end
    always @(spike_out_source_array[995]) begin 
        spike_out_source995 = spike_out_source_array[995];
    end
    always @(spike_out_source_array[996]) begin 
        spike_out_source996 = spike_out_source_array[996];
    end
    always @(spike_out_source_array[997]) begin 
        spike_out_source997 = spike_out_source_array[997];
    end
    always @(spike_out_source_array[998]) begin 
        spike_out_source998 = spike_out_source_array[998];
    end
    always @(spike_out_source_array[999]) begin 
        spike_out_source999 = spike_out_source_array[999];
    end
    always @(spike_out_source_array[1000]) begin 
        spike_out_source1000 = spike_out_source_array[1000];
    end
    always @(spike_out_source_array[1001]) begin 
        spike_out_source1001 = spike_out_source_array[1001];
    end
    always @(spike_out_source_array[1002]) begin 
        spike_out_source1002 = spike_out_source_array[1002];
    end
    always @(spike_out_source_array[1003]) begin 
        spike_out_source1003 = spike_out_source_array[1003];
    end
    always @(spike_out_source_array[1004]) begin 
        spike_out_source1004 = spike_out_source_array[1004];
    end
    always @(spike_out_source_array[1005]) begin 
        spike_out_source1005 = spike_out_source_array[1005];
    end
    always @(spike_out_source_array[1006]) begin 
        spike_out_source1006 = spike_out_source_array[1006];
    end
    always @(spike_out_source_array[1007]) begin 
        spike_out_source1007 = spike_out_source_array[1007];
    end
    always @(spike_out_source_array[1008]) begin 
        spike_out_source1008 = spike_out_source_array[1008];
    end
    always @(spike_out_source_array[1009]) begin 
        spike_out_source1009 = spike_out_source_array[1009];
    end
    always @(spike_out_source_array[1010]) begin 
        spike_out_source1010 = spike_out_source_array[1010];
    end
    always @(spike_out_source_array[1011]) begin 
        spike_out_source1011 = spike_out_source_array[1011];
    end
    always @(spike_out_source_array[1012]) begin 
        spike_out_source1012 = spike_out_source_array[1012];
    end
    always @(spike_out_source_array[1013]) begin 
        spike_out_source1013 = spike_out_source_array[1013];
    end
    always @(spike_out_source_array[1014]) begin 
        spike_out_source1014 = spike_out_source_array[1014];
    end
    always @(spike_out_source_array[1015]) begin 
        spike_out_source1015 = spike_out_source_array[1015];
    end
    always @(spike_out_source_array[1016]) begin 
        spike_out_source1016 = spike_out_source_array[1016];
    end
    always @(spike_out_source_array[1017]) begin 
        spike_out_source1017 = spike_out_source_array[1017];
    end
    always @(spike_out_source_array[1018]) begin 
        spike_out_source1018 = spike_out_source_array[1018];
    end
    always @(spike_out_source_array[1019]) begin 
        spike_out_source1019 = spike_out_source_array[1019];
    end
    always @(spike_out_source_array[1020]) begin 
        spike_out_source1020 = spike_out_source_array[1020];
    end
    always @(spike_out_source_array[1021]) begin 
        spike_out_source1021 = spike_out_source_array[1021];
    end
    always @(spike_out_source_array[1022]) begin 
        spike_out_source1022 = spike_out_source_array[1022];
    end
    always @(spike_out_source_array[1023]) begin 
        spike_out_source1023 = spike_out_source_array[1023];
    end
    reg[18:0] i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21, module network_interface_scaled (
        input wire spike0,
    input wire spike1,    input wire spike2,    input wire spike3,    input wire spike4,    input wire spike5,    input wire spike6,    input wire spike7,    input wire spike8,    input wire spike9,    input wire spike10,    input wire spike11,    input wire spike12,    input wire spike13,    input wire spike14,    input wire spike15,    input wire spike16,    input wire spike17,    input wire spike18,    input wire spike19,    input wire spike20,    input wire spike21,    input wire spike22,    input wire spike23,    input wire spike24,    input wire spike25,    input wire spike26,    input wire spike27,    input wire spike28,    input wire spike29,    input wire spike30,    input wire spike31,    input wire spike32,    input wire spike33,    input wire spike34,    input wire spike35,    input wire spike36,    input wire spike37,    input wire spike38,    input wire spike39,    input wire spike40,    input wire spike41,    input wire spike42,    input wire spike43,    input wire spike44,    input wire spike45,    input wire spike46,    input wire spike47,    input wire spike48,    input wire spike49,    input wire spike50,    input wire spike51,    input wire spike52,    input wire spike53,    input wire spike54,    input wire spike55,    input wire spike56,    input wire spike57,    input wire spike58,    input wire spike59,    input wire spike60,    input wire spike61,    input wire spike62,    input wire spike63,    input wire spike64,    input wire spike65,    input wire spike66,    input wire spike67,    input wire spike68,    input wire spike69,    input wire spike70,    input wire spike71,    input wire spike72,    input wire spike73,    input wire spike74,    input wire spike75,    input wire spike76,    input wire spike77,    input wire spike78,    input wire spike79,    input wire spike80,    input wire spike81,    input wire spike82,    input wire spike83,    input wire spike84,    input wire spike85,    input wire spike86,    input wire spike87,    input wire spike88,    input wire spike89,    input wire spike90,    input wire spike91,    input wire spike92,    input wire spike93,    input wire spike94,    input wire spike95,    input wire spike96,    input wire spike97,    input wire spike98,    input wire spike99,    input wire spike100,
    input wire spike101,    input wire spike102,    input wire spike103,    input wire spike104,    input wire spike105,    input wire spike106,    input wire spike107,    input wire spike108,    input wire spike109,    input wire spike110,    input wire spike111,    input wire spike112,    input wire spike113,    input wire spike114,    input wire spike115,    input wire spike116,    input wire spike117,    input wire spike118,    input wire spike119,    input wire spike120,    input wire spike121,    input wire spike122,    input wire spike123,    input wire spike124,    input wire spike125,    input wire spike126,    input wire spike127,    input wire spike128,    input wire spike129,    input wire spike130,    input wire spike131,    input wire spike132,    input wire spike133,    input wire spike134,    input wire spike135,    input wire spike136,    input wire spike137,    input wire spike138,    input wire spike139,    input wire spike140,    input wire spike141,    input wire spike142,    input wire spike143,    input wire spike144,    input wire spike145,    input wire spike146,    input wire spike147,    input wire spike148,    input wire spike149,    input wire spike150,    input wire spike151,    input wire spike152,    input wire spike153,    input wire spike154,    input wire spike155,    input wire spike156,    input wire spike157,    input wire spike158,    input wire spike159,    input wire spike160,    input wire spike161,    input wire spike162,    input wire spike163,    input wire spike164,    input wire spike165,    input wire spike166,    input wire spike167,    input wire spike168,    input wire spike169,    input wire spike170,    input wire spike171,    input wire spike172,    input wire spike173,    input wire spike174,    input wire spike175,    input wire spike176,    input wire spike177,    input wire spike178,    input wire spike179,    input wire spike180,    input wire spike181,    input wire spike182,    input wire spike183,    input wire spike184,    input wire spike185,    input wire spike186,    input wire spike187,    input wire spike188,    input wire spike189,    input wire spike190,    input wire spike191,    input wire spike192,    input wire spike193,    input wire spike194,    input wire spike195,    input wire spike196,    input wire spike197,    input wire spike198,    input wire spike199,    input wire spike200,
    input wire spike201,    input wire spike202,    input wire spike203,    input wire spike204,    input wire spike205,    input wire spike206,    input wire spike207,    input wire spike208,    input wire spike209,    input wire spike210,    input wire spike211,    input wire spike212,    input wire spike213,    input wire spike214,    input wire spike215,    input wire spike216,    input wire spike217,    input wire spike218,    input wire spike219,    input wire spike220,    input wire spike221,    input wire spike222,    input wire spike223,    input wire spike224,    input wire spike225,    input wire spike226,    input wire spike227,    input wire spike228,    input wire spike229,    input wire spike230,    input wire spike231,    input wire spike232,    input wire spike233,    input wire spike234,    input wire spike235,    input wire spike236,    input wire spike237,    input wire spike238,    input wire spike239,    input wire spike240,    input wire spike241,    input wire spike242,    input wire spike243,    input wire spike244,    input wire spike245,    input wire spike246,    input wire spike247,    input wire spike248,    input wire spike249,    input wire spike250,    input wire spike251,    input wire spike252,    input wire spike253,    input wire spike254,    input wire spike255,    input wire spike256,    input wire spike257,    input wire spike258,    input wire spike259,    input wire spike260,    input wire spike261,    input wire spike262,    input wire spike263,    input wire spike264,    input wire spike265,    input wire spike266,    input wire spike267,    input wire spike268,    input wire spike269,    input wire spike270,    input wire spike271,    input wire spike272,    input wire spike273,    input wire spike274,    input wire spike275,    input wire spike276,    input wire spike277,    input wire spike278,    input wire spike279,    input wire spike280,    input wire spike281,    input wire spike282,    input wire spike283,    input wire spike284,    input wire spike285,    input wire spike286,    input wire spike287,    input wire spike288,    input wire spike289,    input wire spike290,    input wire spike291,    input wire spike292,    input wire spike293,    input wire spike294,    input wire spike295,    input wire spike296,    input wire spike297,    input wire spike298,    input wire spike299,    input wire spike300,
    input wire spike301,    input wire spike302,    input wire spike303,    input wire spike304,    input wire spike305,    input wire spike306,    input wire spike307,    input wire spike308,    input wire spike309,    input wire spike310,    input wire spike311,    input wire spike312,    input wire spike313,    input wire spike314,    input wire spike315,    input wire spike316,    input wire spike317,    input wire spike318,    input wire spike319,    input wire spike320,    input wire spike321,    input wire spike322,    input wire spike323,    input wire spike324,    input wire spike325,    input wire spike326,    input wire spike327,    input wire spike328,    input wire spike329,    input wire spike330,    input wire spike331,    input wire spike332,    input wire spike333,    input wire spike334,    input wire spike335,    input wire spike336,    input wire spike337,    input wire spike338,    input wire spike339,    input wire spike340,    input wire spike341,    input wire spike342,    input wire spike343,    input wire spike344,    input wire spike345,    input wire spike346,    input wire spike347,    input wire spike348,    input wire spike349,    input wire spike350,    input wire spike351,    input wire spike352,    input wire spike353,    input wire spike354,    input wire spike355,    input wire spike356,    input wire spike357,    input wire spike358,    input wire spike359,    input wire spike360,    input wire spike361,    input wire spike362,    input wire spike363,    input wire spike364,    input wire spike365,    input wire spike366,    input wire spike367,    input wire spike368,    input wire spike369,    input wire spike370,    input wire spike371,    input wire spike372,    input wire spike373,    input wire spike374,    input wire spike375,    input wire spike376,    input wire spike377,    input wire spike378,    input wire spike379,    input wire spike380,    input wire spike381,    input wire spike382,    input wire spike383,    input wire spike384,    input wire spike385,    input wire spike386,    input wire spike387,    input wire spike388,    input wire spike389,    input wire spike390,    input wire spike391,    input wire spike392,    input wire spike393,    input wire spike394,    input wire spike395,    input wire spike396,    input wire spike397,    input wire spike398,    input wire spike399,    input wire spike400,
    input wire spike401,    input wire spike402,    input wire spike403,    input wire spike404,    input wire spike405,    input wire spike406,    input wire spike407,    input wire spike408,    input wire spike409,    input wire spike410,    input wire spike411,    input wire spike412,    input wire spike413,    input wire spike414,    input wire spike415,    input wire spike416,    input wire spike417,    input wire spike418,    input wire spike419,    input wire spike420,    input wire spike421,    input wire spike422,    input wire spike423,    input wire spike424,    input wire spike425,    input wire spike426,    input wire spike427,    input wire spike428,    input wire spike429,    input wire spike430,    input wire spike431,    input wire spike432,    input wire spike433,    input wire spike434,    input wire spike435,    input wire spike436,    input wire spike437,    input wire spike438,    input wire spike439,    input wire spike440,    input wire spike441,    input wire spike442,    input wire spike443,    input wire spike444,    input wire spike445,    input wire spike446,    input wire spike447,    input wire spike448,    input wire spike449,    input wire spike450,    input wire spike451,    input wire spike452,    input wire spike453,    input wire spike454,    input wire spike455,    input wire spike456,    input wire spike457,    input wire spike458,    input wire spike459,    input wire spike460,    input wire spike461,    input wire spike462,    input wire spike463,    input wire spike464,    input wire spike465,    input wire spike466,    input wire spike467,    input wire spike468,    input wire spike469,    input wire spike470,    input wire spike471,    input wire spike472,    input wire spike473,    input wire spike474,    input wire spike475,    input wire spike476,    input wire spike477,    input wire spike478,    input wire spike479,    input wire spike480,    input wire spike481,    input wire spike482,    input wire spike483,    input wire spike484,    input wire spike485,    input wire spike486,    input wire spike487,    input wire spike488,    input wire spike489,    input wire spike490,    input wire spike491,    input wire spike492,    input wire spike493,    input wire spike494,    input wire spike495,    input wire spike496,    input wire spike497,    input wire spike498,    input wire spike499,    input wire spike500,
    input wire spike501,    input wire spike502,    input wire spike503,    input wire spike504,    input wire spike505,    input wire spike506,    input wire spike507,    input wire spike508,    input wire spike509,    input wire spike510,    input wire spike511,    input wire spike512,    input wire spike513,    input wire spike514,    input wire spike515,    input wire spike516,    input wire spike517,    input wire spike518,    input wire spike519,    input wire spike520,    input wire spike521,    input wire spike522,    input wire spike523,    input wire spike524,    input wire spike525,    input wire spike526,    input wire spike527,    input wire spike528,    input wire spike529,    input wire spike530,    input wire spike531,    input wire spike532,    input wire spike533,    input wire spike534,    input wire spike535,    input wire spike536,    input wire spike537,    input wire spike538,    input wire spike539,    input wire spike540,    input wire spike541,    input wire spike542,    input wire spike543,    input wire spike544,    input wire spike545,    input wire spike546,    input wire spike547,    input wire spike548,    input wire spike549,    input wire spike550,    input wire spike551,    input wire spike552,    input wire spike553,    input wire spike554,    input wire spike555,    input wire spike556,    input wire spike557,    input wire spike558,    input wire spike559,    input wire spike560,    input wire spike561,    input wire spike562,    input wire spike563,    input wire spike564,    input wire spike565,    input wire spike566,    input wire spike567,    input wire spike568,    input wire spike569,    input wire spike570,    input wire spike571,    input wire spike572,    input wire spike573,    input wire spike574,    input wire spike575,    input wire spike576,    input wire spike577,    input wire spike578,    input wire spike579,    input wire spike580,    input wire spike581,    input wire spike582,    input wire spike583,    input wire spike584,    input wire spike585,    input wire spike586,    input wire spike587,    input wire spike588,    input wire spike589,    input wire spike590,    input wire spike591,    input wire spike592,    input wire spike593,    input wire spike594,    input wire spike595,    input wire spike596,    input wire spike597,    input wire spike598,    input wire spike599,    input wire spike600,
    input wire spike601,    input wire spike602,    input wire spike603,    input wire spike604,    input wire spike605,    input wire spike606,    input wire spike607,    input wire spike608,    input wire spike609,    input wire spike610,    input wire spike611,    input wire spike612,    input wire spike613,    input wire spike614,    input wire spike615,    input wire spike616,    input wire spike617,    input wire spike618,    input wire spike619,    input wire spike620,    input wire spike621,    input wire spike622,    input wire spike623,    input wire spike624,    input wire spike625,    input wire spike626,    input wire spike627,    input wire spike628,    input wire spike629,    input wire spike630,    input wire spike631,    input wire spike632,    input wire spike633,    input wire spike634,    input wire spike635,    input wire spike636,    input wire spike637,    input wire spike638,    input wire spike639,    input wire spike640,    input wire spike641,    input wire spike642,    input wire spike643,    input wire spike644,    input wire spike645,    input wire spike646,    input wire spike647,    input wire spike648,    input wire spike649,    input wire spike650,    input wire spike651,    input wire spike652,    input wire spike653,    input wire spike654,    input wire spike655,    input wire spike656,    input wire spike657,    input wire spike658,    input wire spike659,    input wire spike660,    input wire spike661,    input wire spike662,    input wire spike663,    input wire spike664,    input wire spike665,    input wire spike666,    input wire spike667,    input wire spike668,    input wire spike669,    input wire spike670,    input wire spike671,    input wire spike672,    input wire spike673,    input wire spike674,    input wire spike675,    input wire spike676,    input wire spike677,    input wire spike678,    input wire spike679,    input wire spike680,    input wire spike681,    input wire spike682,    input wire spike683,    input wire spike684,    input wire spike685,    input wire spike686,    input wire spike687,    input wire spike688,    input wire spike689,    input wire spike690,    input wire spike691,    input wire spike692,    input wire spike693,    input wire spike694,    input wire spike695,    input wire spike696,    input wire spike697,    input wire spike698,    input wire spike699,    input wire spike700,
    input wire spike701,    input wire spike702,    input wire spike703,    input wire spike704,    input wire spike705,    input wire spike706,    input wire spike707,    input wire spike708,    input wire spike709,    input wire spike710,    input wire spike711,    input wire spike712,    input wire spike713,    input wire spike714,    input wire spike715,    input wire spike716,    input wire spike717,    input wire spike718,    input wire spike719,    input wire spike720,    input wire spike721,    input wire spike722,    input wire spike723,    input wire spike724,    input wire spike725,    input wire spike726,    input wire spike727,    input wire spike728,    input wire spike729,    input wire spike730,    input wire spike731,    input wire spike732,    input wire spike733,    input wire spike734,    input wire spike735,    input wire spike736,    input wire spike737,    input wire spike738,    input wire spike739,    input wire spike740,    input wire spike741,    input wire spike742,    input wire spike743,    input wire spike744,    input wire spike745,    input wire spike746,    input wire spike747,    input wire spike748,    input wire spike749,    input wire spike750,    input wire spike751,    input wire spike752,    input wire spike753,    input wire spike754,    input wire spike755,    input wire spike756,    input wire spike757,    input wire spike758,    input wire spike759,    input wire spike760,    input wire spike761,    input wire spike762,    input wire spike763,    input wire spike764,    input wire spike765,    input wire spike766,    input wire spike767,    input wire spike768,    input wire spike769,    input wire spike770,    input wire spike771,    input wire spike772,    input wire spike773,    input wire spike774,    input wire spike775,    input wire spike776,    input wire spike777,    input wire spike778,    input wire spike779,    input wire spike780,    input wire spike781,    input wire spike782,    input wire spike783,    input wire spike784,    input wire spike785,    input wire spike786,    input wire spike787,    input wire spike788,    input wire spike789,    input wire spike790,    input wire spike791,    input wire spike792,    input wire spike793,    input wire spike794,    input wire spike795,    input wire spike796,    input wire spike797,    input wire spike798,    input wire spike799,    input wire spike800,
    input wire spike801,    input wire spike802,    input wire spike803,    input wire spike804,    input wire spike805,    input wire spike806,    input wire spike807,    input wire spike808,    input wire spike809,    input wire spike810,    input wire spike811,    input wire spike812,    input wire spike813,    input wire spike814,    input wire spike815,    input wire spike816,    input wire spike817,    input wire spike818,    input wire spike819,    input wire spike820,    input wire spike821,    input wire spike822,    input wire spike823,    input wire spike824,    input wire spike825,    input wire spike826,    input wire spike827,    input wire spike828,    input wire spike829,    input wire spike830,    input wire spike831,    input wire spike832,    input wire spike833,    input wire spike834,    input wire spike835,    input wire spike836,    input wire spike837,    input wire spike838,    input wire spike839,    input wire spike840,    input wire spike841,    input wire spike842,    input wire spike843,    input wire spike844,    input wire spike845,    input wire spike846,    input wire spike847,    input wire spike848,    input wire spike849,    input wire spike850,    input wire spike851,    input wire spike852,    input wire spike853,    input wire spike854,    input wire spike855,    input wire spike856,    input wire spike857,    input wire spike858,    input wire spike859,    input wire spike860,    input wire spike861,    input wire spike862,    input wire spike863,    input wire spike864,    input wire spike865,    input wire spike866,    input wire spike867,    input wire spike868,    input wire spike869,    input wire spike870,    input wire spike871,    input wire spike872,    input wire spike873,    input wire spike874,    input wire spike875,    input wire spike876,    input wire spike877,    input wire spike878,    input wire spike879,    input wire spike880,    input wire spike881,    input wire spike882,    input wire spike883,    input wire spike884,    input wire spike885,    input wire spike886,    input wire spike887,    input wire spike888,    input wire spike889,    input wire spike890,    input wire spike891,    input wire spike892,    input wire spike893,    input wire spike894,    input wire spike895,    input wire spike896,    input wire spike897,    input wire spike898,    input wire spike899,    input wire spike900,
    input wire spike901,    input wire spike902,    input wire spike903,    input wire spike904,    input wire spike905,    input wire spike906,    input wire spike907,    input wire spike908,    input wire spike909,    input wire spike910,    input wire spike911,    input wire spike912,    input wire spike913,    input wire spike914,    input wire spike915,    input wire spike916,    input wire spike917,    input wire spike918,    input wire spike919,    input wire spike920,    input wire spike921,    input wire spike922,    input wire spike923,    input wire spike924,    input wire spike925,    input wire spike926,    input wire spike927,    input wire spike928,    input wire spike929,    input wire spike930,    input wire spike931,    input wire spike932,    input wire spike933,    input wire spike934,    input wire spike935,    input wire spike936,    input wire spike937,    input wire spike938,    input wire spike939,    input wire spike940,    input wire spike941,    input wire spike942,    input wire spike943,    input wire spike944,    input wire spike945,    input wire spike946,    input wire spike947,    input wire spike948,    input wire spike949,    input wire spike950,    input wire spike951,    input wire spike952,    input wire spike953,    input wire spike954,    input wire spike955,    input wire spike956,    input wire spike957,    input wire spike958,    input wire spike959,    input wire spike960,    input wire spike961,    input wire spike962,    input wire spike963,    input wire spike964,    input wire spike965,    input wire spike966,    input wire spike967,    input wire spike968,    input wire spike969,    input wire spike970,    input wire spike971,    input wire spike972,    input wire spike973,    input wire spike974,    input wire spike975,    input wire spike976,    input wire spike977,    input wire spike978,    input wire spike979,    input wire spike980,    input wire spike981,    input wire spike982,    input wire spike983,    input wire spike984,    input wire spike985,    input wire spike986,    input wire spike987,    input wire spike988,    input wire spike989,    input wire spike990,    input wire spike991,    input wire spike992,    input wire spike993,    input wire spike994,    input wire spike995,    input wire spike996,    input wire spike997,    input wire spike998,    input wire spike999,    input wire spike1000,
    input wire spike1001,    input wire spike1002,    input wire spike1003,    input wire spike1004,    input wire spike1005,    input wire spike1006,    input wire spike1007,    input wire spike1008,    input wire spike1009,    input wire spike1010,    input wire spike1011,    input wire spike1012,    input wire spike1013,    input wire spike1014,    input wire spike1015,    input wire spike1016,    input wire spike1017,    input wire spike1018,    input wire spike1019,    input wire spike1020,    input wire spike1021,    input wire spike1022,    input wire spike1023,
output reg[11:0]     spike_out_source0,
    spike_out_source1,    spike_out_source2,    spike_out_source3,    spike_out_source4,    spike_out_source5,    spike_out_source6,    spike_out_source7,    spike_out_source8,    spike_out_source9,    spike_out_source10,    spike_out_source11,    spike_out_source12,    spike_out_source13,    spike_out_source14,    spike_out_source15,    spike_out_source16,    spike_out_source17,    spike_out_source18,    spike_out_source19,    spike_out_source20,    spike_out_source21,    spike_out_source22,    spike_out_source23,    spike_out_source24,    spike_out_source25,    spike_out_source26,    spike_out_source27,    spike_out_source28,    spike_out_source29,    spike_out_source30,    spike_out_source31,    spike_out_source32,    spike_out_source33,    spike_out_source34,    spike_out_source35,    spike_out_source36,    spike_out_source37,    spike_out_source38,    spike_out_source39,    spike_out_source40,    spike_out_source41,    spike_out_source42,    spike_out_source43,    spike_out_source44,    spike_out_source45,    spike_out_source46,    spike_out_source47,    spike_out_source48,    spike_out_source49,    spike_out_source50,    spike_out_source51,    spike_out_source52,    spike_out_source53,    spike_out_source54,    spike_out_source55,    spike_out_source56,    spike_out_source57,    spike_out_source58,    spike_out_source59,    spike_out_source60,    spike_out_source61,    spike_out_source62,    spike_out_source63,    spike_out_source64,    spike_out_source65,    spike_out_source66,    spike_out_source67,    spike_out_source68,    spike_out_source69,    spike_out_source70,    spike_out_source71,    spike_out_source72,    spike_out_source73,    spike_out_source74,    spike_out_source75,    spike_out_source76,    spike_out_source77,    spike_out_source78,    spike_out_source79,    spike_out_source80,    spike_out_source81,    spike_out_source82,    spike_out_source83,    spike_out_source84,    spike_out_source85,    spike_out_source86,    spike_out_source87,    spike_out_source88,    spike_out_source89,    spike_out_source90,    spike_out_source91,    spike_out_source92,    spike_out_source93,    spike_out_source94,    spike_out_source95,    spike_out_source96,    spike_out_source97,    spike_out_source98,    spike_out_source99,    spike_out_source100,
    spike_out_source101,    spike_out_source102,    spike_out_source103,    spike_out_source104,    spike_out_source105,    spike_out_source106,    spike_out_source107,    spike_out_source108,    spike_out_source109,    spike_out_source110,    spike_out_source111,    spike_out_source112,    spike_out_source113,    spike_out_source114,    spike_out_source115,    spike_out_source116,    spike_out_source117,    spike_out_source118,    spike_out_source119,    spike_out_source120,    spike_out_source121,    spike_out_source122,    spike_out_source123,    spike_out_source124,    spike_out_source125,    spike_out_source126,    spike_out_source127,    spike_out_source128,    spike_out_source129,    spike_out_source130,    spike_out_source131,    spike_out_source132,    spike_out_source133,    spike_out_source134,    spike_out_source135,    spike_out_source136,    spike_out_source137,    spike_out_source138,    spike_out_source139,    spike_out_source140,    spike_out_source141,    spike_out_source142,    spike_out_source143,    spike_out_source144,    spike_out_source145,    spike_out_source146,    spike_out_source147,    spike_out_source148,    spike_out_source149,    spike_out_source150,    spike_out_source151,    spike_out_source152,    spike_out_source153,    spike_out_source154,    spike_out_source155,    spike_out_source156,    spike_out_source157,    spike_out_source158,    spike_out_source159,    spike_out_source160,    spike_out_source161,    spike_out_source162,    spike_out_source163,    spike_out_source164,    spike_out_source165,    spike_out_source166,    spike_out_source167,    spike_out_source168,    spike_out_source169,    spike_out_source170,    spike_out_source171,    spike_out_source172,    spike_out_source173,    spike_out_source174,    spike_out_source175,    spike_out_source176,    spike_out_source177,    spike_out_source178,    spike_out_source179,    spike_out_source180,    spike_out_source181,    spike_out_source182,    spike_out_source183,    spike_out_source184,    spike_out_source185,    spike_out_source186,    spike_out_source187,    spike_out_source188,    spike_out_source189,    spike_out_source190,    spike_out_source191,    spike_out_source192,    spike_out_source193,    spike_out_source194,    spike_out_source195,    spike_out_source196,    spike_out_source197,    spike_out_source198,    spike_out_source199,    spike_out_source200,
    spike_out_source201,    spike_out_source202,    spike_out_source203,    spike_out_source204,    spike_out_source205,    spike_out_source206,    spike_out_source207,    spike_out_source208,    spike_out_source209,    spike_out_source210,    spike_out_source211,    spike_out_source212,    spike_out_source213,    spike_out_source214,    spike_out_source215,    spike_out_source216,    spike_out_source217,    spike_out_source218,    spike_out_source219,    spike_out_source220,    spike_out_source221,    spike_out_source222,    spike_out_source223,    spike_out_source224,    spike_out_source225,    spike_out_source226,    spike_out_source227,    spike_out_source228,    spike_out_source229,    spike_out_source230,    spike_out_source231,    spike_out_source232,    spike_out_source233,    spike_out_source234,    spike_out_source235,    spike_out_source236,    spike_out_source237,    spike_out_source238,    spike_out_source239,    spike_out_source240,    spike_out_source241,    spike_out_source242,    spike_out_source243,    spike_out_source244,    spike_out_source245,    spike_out_source246,    spike_out_source247,    spike_out_source248,    spike_out_source249,    spike_out_source250,    spike_out_source251,    spike_out_source252,    spike_out_source253,    spike_out_source254,    spike_out_source255,    spike_out_source256,    spike_out_source257,    spike_out_source258,    spike_out_source259,    spike_out_source260,    spike_out_source261,    spike_out_source262,    spike_out_source263,    spike_out_source264,    spike_out_source265,    spike_out_source266,    spike_out_source267,    spike_out_source268,    spike_out_source269,    spike_out_source270,    spike_out_source271,    spike_out_source272,    spike_out_source273,    spike_out_source274,    spike_out_source275,    spike_out_source276,    spike_out_source277,    spike_out_source278,    spike_out_source279,    spike_out_source280,    spike_out_source281,    spike_out_source282,    spike_out_source283,    spike_out_source284,    spike_out_source285,    spike_out_source286,    spike_out_source287,    spike_out_source288,    spike_out_source289,    spike_out_source290,    spike_out_source291,    spike_out_source292,    spike_out_source293,    spike_out_source294,    spike_out_source295,    spike_out_source296,    spike_out_source297,    spike_out_source298,    spike_out_source299,    spike_out_source300,
    spike_out_source301,    spike_out_source302,    spike_out_source303,    spike_out_source304,    spike_out_source305,    spike_out_source306,    spike_out_source307,    spike_out_source308,    spike_out_source309,    spike_out_source310,    spike_out_source311,    spike_out_source312,    spike_out_source313,    spike_out_source314,    spike_out_source315,    spike_out_source316,    spike_out_source317,    spike_out_source318,    spike_out_source319,    spike_out_source320,    spike_out_source321,    spike_out_source322,    spike_out_source323,    spike_out_source324,    spike_out_source325,    spike_out_source326,    spike_out_source327,    spike_out_source328,    spike_out_source329,    spike_out_source330,    spike_out_source331,    spike_out_source332,    spike_out_source333,    spike_out_source334,    spike_out_source335,    spike_out_source336,    spike_out_source337,    spike_out_source338,    spike_out_source339,    spike_out_source340,    spike_out_source341,    spike_out_source342,    spike_out_source343,    spike_out_source344,    spike_out_source345,    spike_out_source346,    spike_out_source347,    spike_out_source348,    spike_out_source349,    spike_out_source350,    spike_out_source351,    spike_out_source352,    spike_out_source353,    spike_out_source354,    spike_out_source355,    spike_out_source356,    spike_out_source357,    spike_out_source358,    spike_out_source359,    spike_out_source360,    spike_out_source361,    spike_out_source362,    spike_out_source363,    spike_out_source364,    spike_out_source365,    spike_out_source366,    spike_out_source367,    spike_out_source368,    spike_out_source369,    spike_out_source370,    spike_out_source371,    spike_out_source372,    spike_out_source373,    spike_out_source374,    spike_out_source375,    spike_out_source376,    spike_out_source377,    spike_out_source378,    spike_out_source379,    spike_out_source380,    spike_out_source381,    spike_out_source382,    spike_out_source383,    spike_out_source384,    spike_out_source385,    spike_out_source386,    spike_out_source387,    spike_out_source388,    spike_out_source389,    spike_out_source390,    spike_out_source391,    spike_out_source392,    spike_out_source393,    spike_out_source394,    spike_out_source395,    spike_out_source396,    spike_out_source397,    spike_out_source398,    spike_out_source399,    spike_out_source400,
    spike_out_source401,    spike_out_source402,    spike_out_source403,    spike_out_source404,    spike_out_source405,    spike_out_source406,    spike_out_source407,    spike_out_source408,    spike_out_source409,    spike_out_source410,    spike_out_source411,    spike_out_source412,    spike_out_source413,    spike_out_source414,    spike_out_source415,    spike_out_source416,    spike_out_source417,    spike_out_source418,    spike_out_source419,    spike_out_source420,    spike_out_source421,    spike_out_source422,    spike_out_source423,    spike_out_source424,    spike_out_source425,    spike_out_source426,    spike_out_source427,    spike_out_source428,    spike_out_source429,    spike_out_source430,    spike_out_source431,    spike_out_source432,    spike_out_source433,    spike_out_source434,    spike_out_source435,    spike_out_source436,    spike_out_source437,    spike_out_source438,    spike_out_source439,    spike_out_source440,    spike_out_source441,    spike_out_source442,    spike_out_source443,    spike_out_source444,    spike_out_source445,    spike_out_source446,    spike_out_source447,    spike_out_source448,    spike_out_source449,    spike_out_source450,    spike_out_source451,    spike_out_source452,    spike_out_source453,    spike_out_source454,    spike_out_source455,    spike_out_source456,    spike_out_source457,    spike_out_source458,    spike_out_source459,    spike_out_source460,    spike_out_source461,    spike_out_source462,    spike_out_source463,    spike_out_source464,    spike_out_source465,    spike_out_source466,    spike_out_source467,    spike_out_source468,    spike_out_source469,    spike_out_source470,    spike_out_source471,    spike_out_source472,    spike_out_source473,    spike_out_source474,    spike_out_source475,    spike_out_source476,    spike_out_source477,    spike_out_source478,    spike_out_source479,    spike_out_source480,    spike_out_source481,    spike_out_source482,    spike_out_source483,    spike_out_source484,    spike_out_source485,    spike_out_source486,    spike_out_source487,    spike_out_source488,    spike_out_source489,    spike_out_source490,    spike_out_source491,    spike_out_source492,    spike_out_source493,    spike_out_source494,    spike_out_source495,    spike_out_source496,    spike_out_source497,    spike_out_source498,    spike_out_source499,    spike_out_source500,
    spike_out_source501,    spike_out_source502,    spike_out_source503,    spike_out_source504,    spike_out_source505,    spike_out_source506,    spike_out_source507,    spike_out_source508,    spike_out_source509,    spike_out_source510,    spike_out_source511,    spike_out_source512,    spike_out_source513,    spike_out_source514,    spike_out_source515,    spike_out_source516,    spike_out_source517,    spike_out_source518,    spike_out_source519,    spike_out_source520,    spike_out_source521,    spike_out_source522,    spike_out_source523,    spike_out_source524,    spike_out_source525,    spike_out_source526,    spike_out_source527,    spike_out_source528,    spike_out_source529,    spike_out_source530,    spike_out_source531,    spike_out_source532,    spike_out_source533,    spike_out_source534,    spike_out_source535,    spike_out_source536,    spike_out_source537,    spike_out_source538,    spike_out_source539,    spike_out_source540,    spike_out_source541,    spike_out_source542,    spike_out_source543,    spike_out_source544,    spike_out_source545,    spike_out_source546,    spike_out_source547,    spike_out_source548,    spike_out_source549,    spike_out_source550,    spike_out_source551,    spike_out_source552,    spike_out_source553,    spike_out_source554,    spike_out_source555,    spike_out_source556,    spike_out_source557,    spike_out_source558,    spike_out_source559,    spike_out_source560,    spike_out_source561,    spike_out_source562,    spike_out_source563,    spike_out_source564,    spike_out_source565,    spike_out_source566,    spike_out_source567,    spike_out_source568,    spike_out_source569,    spike_out_source570,    spike_out_source571,    spike_out_source572,    spike_out_source573,    spike_out_source574,    spike_out_source575,    spike_out_source576,    spike_out_source577,    spike_out_source578,    spike_out_source579,    spike_out_source580,    spike_out_source581,    spike_out_source582,    spike_out_source583,    spike_out_source584,    spike_out_source585,    spike_out_source586,    spike_out_source587,    spike_out_source588,    spike_out_source589,    spike_out_source590,    spike_out_source591,    spike_out_source592,    spike_out_source593,    spike_out_source594,    spike_out_source595,    spike_out_source596,    spike_out_source597,    spike_out_source598,    spike_out_source599,    spike_out_source600,
    spike_out_source601,    spike_out_source602,    spike_out_source603,    spike_out_source604,    spike_out_source605,    spike_out_source606,    spike_out_source607,    spike_out_source608,    spike_out_source609,    spike_out_source610,    spike_out_source611,    spike_out_source612,    spike_out_source613,    spike_out_source614,    spike_out_source615,    spike_out_source616,    spike_out_source617,    spike_out_source618,    spike_out_source619,    spike_out_source620,    spike_out_source621,    spike_out_source622,    spike_out_source623,    spike_out_source624,    spike_out_source625,    spike_out_source626,    spike_out_source627,    spike_out_source628,    spike_out_source629,    spike_out_source630,    spike_out_source631,    spike_out_source632,    spike_out_source633,    spike_out_source634,    spike_out_source635,    spike_out_source636,    spike_out_source637,    spike_out_source638,    spike_out_source639,    spike_out_source640,    spike_out_source641,    spike_out_source642,    spike_out_source643,    spike_out_source644,    spike_out_source645,    spike_out_source646,    spike_out_source647,    spike_out_source648,    spike_out_source649,    spike_out_source650,    spike_out_source651,    spike_out_source652,    spike_out_source653,    spike_out_source654,    spike_out_source655,    spike_out_source656,    spike_out_source657,    spike_out_source658,    spike_out_source659,    spike_out_source660,    spike_out_source661,    spike_out_source662,    spike_out_source663,    spike_out_source664,    spike_out_source665,    spike_out_source666,    spike_out_source667,    spike_out_source668,    spike_out_source669,    spike_out_source670,    spike_out_source671,    spike_out_source672,    spike_out_source673,    spike_out_source674,    spike_out_source675,    spike_out_source676,    spike_out_source677,    spike_out_source678,    spike_out_source679,    spike_out_source680,    spike_out_source681,    spike_out_source682,    spike_out_source683,    spike_out_source684,    spike_out_source685,    spike_out_source686,    spike_out_source687,    spike_out_source688,    spike_out_source689,    spike_out_source690,    spike_out_source691,    spike_out_source692,    spike_out_source693,    spike_out_source694,    spike_out_source695,    spike_out_source696,    spike_out_source697,    spike_out_source698,    spike_out_source699,    spike_out_source700,
    spike_out_source701,    spike_out_source702,    spike_out_source703,    spike_out_source704,    spike_out_source705,    spike_out_source706,    spike_out_source707,    spike_out_source708,    spike_out_source709,    spike_out_source710,    spike_out_source711,    spike_out_source712,    spike_out_source713,    spike_out_source714,    spike_out_source715,    spike_out_source716,    spike_out_source717,    spike_out_source718,    spike_out_source719,    spike_out_source720,    spike_out_source721,    spike_out_source722,    spike_out_source723,    spike_out_source724,    spike_out_source725,    spike_out_source726,    spike_out_source727,    spike_out_source728,    spike_out_source729,    spike_out_source730,    spike_out_source731,    spike_out_source732,    spike_out_source733,    spike_out_source734,    spike_out_source735,    spike_out_source736,    spike_out_source737,    spike_out_source738,    spike_out_source739,    spike_out_source740,    spike_out_source741,    spike_out_source742,    spike_out_source743,    spike_out_source744,    spike_out_source745,    spike_out_source746,    spike_out_source747,    spike_out_source748,    spike_out_source749,    spike_out_source750,    spike_out_source751,    spike_out_source752,    spike_out_source753,    spike_out_source754,    spike_out_source755,    spike_out_source756,    spike_out_source757,    spike_out_source758,    spike_out_source759,    spike_out_source760,    spike_out_source761,    spike_out_source762,    spike_out_source763,    spike_out_source764,    spike_out_source765,    spike_out_source766,    spike_out_source767,    spike_out_source768,    spike_out_source769,    spike_out_source770,    spike_out_source771,    spike_out_source772,    spike_out_source773,    spike_out_source774,    spike_out_source775,    spike_out_source776,    spike_out_source777,    spike_out_source778,    spike_out_source779,    spike_out_source780,    spike_out_source781,    spike_out_source782,    spike_out_source783,    spike_out_source784,    spike_out_source785,    spike_out_source786,    spike_out_source787,    spike_out_source788,    spike_out_source789,    spike_out_source790,    spike_out_source791,    spike_out_source792,    spike_out_source793,    spike_out_source794,    spike_out_source795,    spike_out_source796,    spike_out_source797,    spike_out_source798,    spike_out_source799,    spike_out_source800,
    spike_out_source801,    spike_out_source802,    spike_out_source803,    spike_out_source804,    spike_out_source805,    spike_out_source806,    spike_out_source807,    spike_out_source808,    spike_out_source809,    spike_out_source810,    spike_out_source811,    spike_out_source812,    spike_out_source813,    spike_out_source814,    spike_out_source815,    spike_out_source816,    spike_out_source817,    spike_out_source818,    spike_out_source819,    spike_out_source820,    spike_out_source821,    spike_out_source822,    spike_out_source823,    spike_out_source824,    spike_out_source825,    spike_out_source826,    spike_out_source827,    spike_out_source828,    spike_out_source829,    spike_out_source830,    spike_out_source831,    spike_out_source832,    spike_out_source833,    spike_out_source834,    spike_out_source835,    spike_out_source836,    spike_out_source837,    spike_out_source838,    spike_out_source839,    spike_out_source840,    spike_out_source841,    spike_out_source842,    spike_out_source843,    spike_out_source844,    spike_out_source845,    spike_out_source846,    spike_out_source847,    spike_out_source848,    spike_out_source849,    spike_out_source850,    spike_out_source851,    spike_out_source852,    spike_out_source853,    spike_out_source854,    spike_out_source855,    spike_out_source856,    spike_out_source857,    spike_out_source858,    spike_out_source859,    spike_out_source860,    spike_out_source861,    spike_out_source862,    spike_out_source863,    spike_out_source864,    spike_out_source865,    spike_out_source866,    spike_out_source867,    spike_out_source868,    spike_out_source869,    spike_out_source870,    spike_out_source871,    spike_out_source872,    spike_out_source873,    spike_out_source874,    spike_out_source875,    spike_out_source876,    spike_out_source877,    spike_out_source878,    spike_out_source879,    spike_out_source880,    spike_out_source881,    spike_out_source882,    spike_out_source883,    spike_out_source884,    spike_out_source885,    spike_out_source886,    spike_out_source887,    spike_out_source888,    spike_out_source889,    spike_out_source890,    spike_out_source891,    spike_out_source892,    spike_out_source893,    spike_out_source894,    spike_out_source895,    spike_out_source896,    spike_out_source897,    spike_out_source898,    spike_out_source899,    spike_out_source900,
    spike_out_source901,    spike_out_source902,    spike_out_source903,    spike_out_source904,    spike_out_source905,    spike_out_source906,    spike_out_source907,    spike_out_source908,    spike_out_source909,    spike_out_source910,    spike_out_source911,    spike_out_source912,    spike_out_source913,    spike_out_source914,    spike_out_source915,    spike_out_source916,    spike_out_source917,    spike_out_source918,    spike_out_source919,    spike_out_source920,    spike_out_source921,    spike_out_source922,    spike_out_source923,    spike_out_source924,    spike_out_source925,    spike_out_source926,    spike_out_source927,    spike_out_source928,    spike_out_source929,    spike_out_source930,    spike_out_source931,    spike_out_source932,    spike_out_source933,    spike_out_source934,    spike_out_source935,    spike_out_source936,    spike_out_source937,    spike_out_source938,    spike_out_source939,    spike_out_source940,    spike_out_source941,    spike_out_source942,    spike_out_source943,    spike_out_source944,    spike_out_source945,    spike_out_source946,    spike_out_source947,    spike_out_source948,    spike_out_source949,    spike_out_source950,    spike_out_source951,    spike_out_source952,    spike_out_source953,    spike_out_source954,    spike_out_source955,    spike_out_source956,    spike_out_source957,    spike_out_source958,    spike_out_source959,    spike_out_source960,    spike_out_source961,    spike_out_source962,    spike_out_source963,    spike_out_source964,    spike_out_source965,    spike_out_source966,    spike_out_source967,    spike_out_source968,    spike_out_source969,    spike_out_source970,    spike_out_source971,    spike_out_source972,    spike_out_source973,    spike_out_source974,    spike_out_source975,    spike_out_source976,    spike_out_source977,    spike_out_source978,    spike_out_source979,    spike_out_source980,    spike_out_source981,    spike_out_source982,    spike_out_source983,    spike_out_source984,    spike_out_source985,    spike_out_source986,    spike_out_source987,    spike_out_source988,    spike_out_source989,    spike_out_source990,    spike_out_source991,    spike_out_source992,    spike_out_source993,    spike_out_source994,    spike_out_source995,    spike_out_source996,    spike_out_source997,    spike_out_source998,    spike_out_source999,    spike_out_source1000,
    spike_out_source1001,    spike_out_source1002,    spike_out_source1003,    spike_out_source1004,    spike_out_source1005,    spike_out_source1006,    spike_out_source1007,    spike_out_source1008,    spike_out_source1009,    spike_out_source1010,    spike_out_source1011,    spike_out_source1012,    spike_out_source1013,    spike_out_source1014,    spike_out_source1015,    spike_out_source1016,    spike_out_source1017,    spike_out_source1018,    spike_out_source1019,    spike_out_source1020,    spike_out_source1021,    spike_out_source1022,    spike_out_source1023,
    output wire output
);

    parameter number_of_neurons= 1024;
    reg spike_register[0:number_of_neurons-1];
    always @(clear, lock1, spike0, spike1, spike2, spike3, spike4, spike5, spike6, spike7, spike8, spike9, spike10, spike11, spike12, spike13, spike14, spike15, spike16, spike17, spike18, spike19, spike20, spike21, spike22, spike23, spike24, spike25, spike26, spike27, spike28, spike29, spike30, spike31, spike32, spike33, spike34, spike35, spike36, spike37, spike38, spike39, spike40, spike41, spike42, spike43, spike44, spike45, spike46, spike47, spike48, spike49) begin
        spike_register[0] = spike0;

        spike_register[1] = spike1;        spike_register[2] = spike2;        spike_register[3] = spike3;        spike_register[4] = spike4;        spike_register[5] = spike5;        spike_register[6] = spike6;        spike_register[7] = spike7;        spike_register[8] = spike8;        spike_register[9] = spike9;        spike_register[10] = spike10;        spike_register[11] = spike11;        spike_register[12] = spike12;        spike_register[13] = spike13;        spike_register[14] = spike14;        spike_register[15] = spike15;        spike_register[16] = spike16;        spike_register[17] = spike17;        spike_register[18] = spike18;        spike_register[19] = spike19;        spike_register[20] = spike20;        spike_register[21] = spike21;        spike_register[22] = spike22;        spike_register[23] = spike23;        spike_register[24] = spike24;        spike_register[25] = spike25;        spike_register[26] = spike26;        spike_register[27] = spike27;        spike_register[28] = spike28;        spike_register[29] = spike29;        spike_register[30] = spike30;        spike_register[31] = spike31;        spike_register[32] = spike32;        spike_register[33] = spike33;        spike_register[34] = spike34;        spike_register[35] = spike35;        spike_register[36] = spike36;        spike_register[37] = spike37;        spike_register[38] = spike38;        spike_register[39] = spike39;        spike_register[40] = spike40;        spike_register[41] = spike41;        spike_register[42] = spike42;        spike_register[43] = spike43;        spike_register[44] = spike44;        spike_register[45] = spike45;        spike_register[46] = spike46;        spike_register[47] = spike47;        spike_register[48] = spike48;        spike_register[49] = spike49;
        #0.5
        if(clear == 1'b0) begin
            for(i1 = 0; i1 <=49; i1= i1+1) begin
                if(spike_register[i1] == 1 && lock1 == 0) begin
                    lock1 = 1;
                    for(j1 = connection_pointer[i1]; j1 < connection_pointer[i1+1]; j1= j1+1) begin
                        packet1 = #0.1 {neuron_addresses[i1], downstream_connections[j1]};
                    end
                    spike_register[i1] = 0;
                    lock1 = 0;
                end
            end
        end

    end
    always @(clear, lock2, spike50, spike51, spike52, spike53, spike54, spike55, spike56, spike57, spike58, spike59, spike60, spike61, spike62, spike63, spike64, spike65, spike66, spike67, spike68, spike69, spike70, spike71, spike72, spike73, spike74, spike75, spike76, spike77, spike78, spike79, spike80, spike81, spike82, spike83, spike84, spike85, spike86, spike87, spike88, spike89, spike90, spike91, spike92, spike93, spike94, spike95, spike96, spike97, spike98, spike99) begin
        spike_register[50] = spike50;        spike_register[51] = spike51;        spike_register[52] = spike52;        spike_register[53] = spike53;        spike_register[54] = spike54;        spike_register[55] = spike55;        spike_register[56] = spike56;        spike_register[57] = spike57;        spike_register[58] = spike58;        spike_register[59] = spike59;        spike_register[60] = spike60;        spike_register[61] = spike61;        spike_register[62] = spike62;        spike_register[63] = spike63;        spike_register[64] = spike64;        spike_register[65] = spike65;        spike_register[66] = spike66;        spike_register[67] = spike67;        spike_register[68] = spike68;        spike_register[69] = spike69;        spike_register[70] = spike70;        spike_register[71] = spike71;        spike_register[72] = spike72;        spike_register[73] = spike73;        spike_register[74] = spike74;        spike_register[75] = spike75;        spike_register[76] = spike76;        spike_register[77] = spike77;        spike_register[78] = spike78;        spike_register[79] = spike79;        spike_register[80] = spike80;        spike_register[81] = spike81;        spike_register[82] = spike82;        spike_register[83] = spike83;        spike_register[84] = spike84;        spike_register[85] = spike85;        spike_register[86] = spike86;        spike_register[87] = spike87;        spike_register[88] = spike88;        spike_register[89] = spike89;        spike_register[90] = spike90;        spike_register[91] = spike91;        spike_register[92] = spike92;        spike_register[93] = spike93;        spike_register[94] = spike94;        spike_register[95] = spike95;        spike_register[96] = spike96;        spike_register[97] = spike97;        spike_register[98] = spike98;        spike_register[99] = spike99;
        #0.5
        if(clear == 1'b0) begin
            for(i2 = 50; i2 <=99; i2= i2+1) begin
                if(spike_register[i2] == 1 && lock2 == 0) begin
                    lock2 = 1;
                    for(j2 = connection_pointer[i2]; j2 < connection_pointer[i2+1]; j2= j2+1) begin
                        packet2 = #0.1 {neuron_addresses[i2], downstream_connections[j2]};
                    end
                    spike_register[i2] = 0;
                    lock2 = 0;
                end
            end
        end

    end
    always @(clear, lock3, spike100, spike101, spike102, spike103, spike104, spike105, spike106, spike107, spike108, spike109, spike110, spike111, spike112, spike113, spike114, spike115, spike116, spike117, spike118, spike119, spike120, spike121, spike122, spike123, spike124, spike125, spike126, spike127, spike128, spike129, spike130, spike131, spike132, spike133, spike134, spike135, spike136, spike137, spike138, spike139, spike140, spike141, spike142, spike143, spike144, spike145, spike146, spike147, spike148, spike149) begin
        spike_register[100] = spike100;

        spike_register[101] = spike101;        spike_register[102] = spike102;        spike_register[103] = spike103;        spike_register[104] = spike104;        spike_register[105] = spike105;        spike_register[106] = spike106;        spike_register[107] = spike107;        spike_register[108] = spike108;        spike_register[109] = spike109;        spike_register[110] = spike110;        spike_register[111] = spike111;        spike_register[112] = spike112;        spike_register[113] = spike113;        spike_register[114] = spike114;        spike_register[115] = spike115;        spike_register[116] = spike116;        spike_register[117] = spike117;        spike_register[118] = spike118;        spike_register[119] = spike119;        spike_register[120] = spike120;        spike_register[121] = spike121;        spike_register[122] = spike122;        spike_register[123] = spike123;        spike_register[124] = spike124;        spike_register[125] = spike125;        spike_register[126] = spike126;        spike_register[127] = spike127;        spike_register[128] = spike128;        spike_register[129] = spike129;        spike_register[130] = spike130;        spike_register[131] = spike131;        spike_register[132] = spike132;        spike_register[133] = spike133;        spike_register[134] = spike134;        spike_register[135] = spike135;        spike_register[136] = spike136;        spike_register[137] = spike137;        spike_register[138] = spike138;        spike_register[139] = spike139;        spike_register[140] = spike140;        spike_register[141] = spike141;        spike_register[142] = spike142;        spike_register[143] = spike143;        spike_register[144] = spike144;        spike_register[145] = spike145;        spike_register[146] = spike146;        spike_register[147] = spike147;        spike_register[148] = spike148;        spike_register[149] = spike149;
        #0.5
        if(clear == 1'b0) begin
            for(i3 = 100; i3 <=149; i3= i3+1) begin
                if(spike_register[i3] == 1 && lock3 == 0) begin
                    lock3 = 1;
                    for(j3 = connection_pointer[i3]; j3 < connection_pointer[i3+1]; j3= j3+1) begin
                        packet3 = #0.1 {neuron_addresses[i3], downstream_connections[j3]};
                    end
                    spike_register[i3] = 0;
                    lock3 = 0;
                end
            end
        end

    end
    always @(clear, lock4, spike150, spike151, spike152, spike153, spike154, spike155, spike156, spike157, spike158, spike159, spike160, spike161, spike162, spike163, spike164, spike165, spike166, spike167, spike168, spike169, spike170, spike171, spike172, spike173, spike174, spike175, spike176, spike177, spike178, spike179, spike180, spike181, spike182, spike183, spike184, spike185, spike186, spike187, spike188, spike189, spike190, spike191, spike192, spike193, spike194, spike195, spike196, spike197, spike198, spike199) begin
        spike_register[150] = spike150;        spike_register[151] = spike151;        spike_register[152] = spike152;        spike_register[153] = spike153;        spike_register[154] = spike154;        spike_register[155] = spike155;        spike_register[156] = spike156;        spike_register[157] = spike157;        spike_register[158] = spike158;        spike_register[159] = spike159;        spike_register[160] = spike160;        spike_register[161] = spike161;        spike_register[162] = spike162;        spike_register[163] = spike163;        spike_register[164] = spike164;        spike_register[165] = spike165;        spike_register[166] = spike166;        spike_register[167] = spike167;        spike_register[168] = spike168;        spike_register[169] = spike169;        spike_register[170] = spike170;        spike_register[171] = spike171;        spike_register[172] = spike172;        spike_register[173] = spike173;        spike_register[174] = spike174;        spike_register[175] = spike175;        spike_register[176] = spike176;        spike_register[177] = spike177;        spike_register[178] = spike178;        spike_register[179] = spike179;        spike_register[180] = spike180;        spike_register[181] = spike181;        spike_register[182] = spike182;        spike_register[183] = spike183;        spike_register[184] = spike184;        spike_register[185] = spike185;        spike_register[186] = spike186;        spike_register[187] = spike187;        spike_register[188] = spike188;        spike_register[189] = spike189;        spike_register[190] = spike190;        spike_register[191] = spike191;        spike_register[192] = spike192;        spike_register[193] = spike193;        spike_register[194] = spike194;        spike_register[195] = spike195;        spike_register[196] = spike196;        spike_register[197] = spike197;        spike_register[198] = spike198;        spike_register[199] = spike199;
        #0.5
        if(clear == 1'b0) begin
            for(i4 = 150; i4 <=199; i4= i4+1) begin
                if(spike_register[i4] == 1 && lock4 == 0) begin
                    lock4 = 1;
                    for(j4 = connection_pointer[i4]; j4 < connection_pointer[i4+1]; j4= j4+1) begin
                        packet4 = #0.1 {neuron_addresses[i4], downstream_connections[j4]};
                    end
                    spike_register[i4] = 0;
                    lock4 = 0;
                end
            end
        end

    end
    always @(clear, lock5, spike200, spike201, spike202, spike203, spike204, spike205, spike206, spike207, spike208, spike209, spike210, spike211, spike212, spike213, spike214, spike215, spike216, spike217, spike218, spike219, spike220, spike221, spike222, spike223, spike224, spike225, spike226, spike227, spike228, spike229, spike230, spike231, spike232, spike233, spike234, spike235, spike236, spike237, spike238, spike239, spike240, spike241, spike242, spike243, spike244, spike245, spike246, spike247, spike248, spike249) begin
        spike_register[200] = spike200;

        spike_register[201] = spike201;        spike_register[202] = spike202;        spike_register[203] = spike203;        spike_register[204] = spike204;        spike_register[205] = spike205;        spike_register[206] = spike206;        spike_register[207] = spike207;        spike_register[208] = spike208;        spike_register[209] = spike209;        spike_register[210] = spike210;        spike_register[211] = spike211;        spike_register[212] = spike212;        spike_register[213] = spike213;        spike_register[214] = spike214;        spike_register[215] = spike215;        spike_register[216] = spike216;        spike_register[217] = spike217;        spike_register[218] = spike218;        spike_register[219] = spike219;        spike_register[220] = spike220;        spike_register[221] = spike221;        spike_register[222] = spike222;        spike_register[223] = spike223;        spike_register[224] = spike224;        spike_register[225] = spike225;        spike_register[226] = spike226;        spike_register[227] = spike227;        spike_register[228] = spike228;        spike_register[229] = spike229;        spike_register[230] = spike230;        spike_register[231] = spike231;        spike_register[232] = spike232;        spike_register[233] = spike233;        spike_register[234] = spike234;        spike_register[235] = spike235;        spike_register[236] = spike236;        spike_register[237] = spike237;        spike_register[238] = spike238;        spike_register[239] = spike239;        spike_register[240] = spike240;        spike_register[241] = spike241;        spike_register[242] = spike242;        spike_register[243] = spike243;        spike_register[244] = spike244;        spike_register[245] = spike245;        spike_register[246] = spike246;        spike_register[247] = spike247;        spike_register[248] = spike248;        spike_register[249] = spike249;
        #0.5
        if(clear == 1'b0) begin
            for(i5 = 200; i5 <=249; i5= i5+1) begin
                if(spike_register[i5] == 1 && lock5 == 0) begin
                    lock5 = 1;
                    for(j5 = connection_pointer[i5]; j5 < connection_pointer[i5+1]; j5= j5+1) begin
                        packet5 = #0.1 {neuron_addresses[i5], downstream_connections[j5]};
                    end
                    spike_register[i5] = 0;
                    lock5 = 0;
                end
            end
        end

    end
    always @(clear, lock6, spike250, spike251, spike252, spike253, spike254, spike255, spike256, spike257, spike258, spike259, spike260, spike261, spike262, spike263, spike264, spike265, spike266, spike267, spike268, spike269, spike270, spike271, spike272, spike273, spike274, spike275, spike276, spike277, spike278, spike279, spike280, spike281, spike282, spike283, spike284, spike285, spike286, spike287, spike288, spike289, spike290, spike291, spike292, spike293, spike294, spike295, spike296, spike297, spike298, spike299) begin
        spike_register[250] = spike250;        spike_register[251] = spike251;        spike_register[252] = spike252;        spike_register[253] = spike253;        spike_register[254] = spike254;        spike_register[255] = spike255;        spike_register[256] = spike256;        spike_register[257] = spike257;        spike_register[258] = spike258;        spike_register[259] = spike259;        spike_register[260] = spike260;        spike_register[261] = spike261;        spike_register[262] = spike262;        spike_register[263] = spike263;        spike_register[264] = spike264;        spike_register[265] = spike265;        spike_register[266] = spike266;        spike_register[267] = spike267;        spike_register[268] = spike268;        spike_register[269] = spike269;        spike_register[270] = spike270;        spike_register[271] = spike271;        spike_register[272] = spike272;        spike_register[273] = spike273;        spike_register[274] = spike274;        spike_register[275] = spike275;        spike_register[276] = spike276;        spike_register[277] = spike277;        spike_register[278] = spike278;        spike_register[279] = spike279;        spike_register[280] = spike280;        spike_register[281] = spike281;        spike_register[282] = spike282;        spike_register[283] = spike283;        spike_register[284] = spike284;        spike_register[285] = spike285;        spike_register[286] = spike286;        spike_register[287] = spike287;        spike_register[288] = spike288;        spike_register[289] = spike289;        spike_register[290] = spike290;        spike_register[291] = spike291;        spike_register[292] = spike292;        spike_register[293] = spike293;        spike_register[294] = spike294;        spike_register[295] = spike295;        spike_register[296] = spike296;        spike_register[297] = spike297;        spike_register[298] = spike298;        spike_register[299] = spike299;
        #0.5
        if(clear == 1'b0) begin
            for(i6 = 250; i6 <=299; i6= i6+1) begin
                if(spike_register[i6] == 1 && lock6 == 0) begin
                    lock6 = 1;
                    for(j6 = connection_pointer[i6]; j6 < connection_pointer[i6+1]; j6= j6+1) begin
                        packet6 = #0.1 {neuron_addresses[i6], downstream_connections[j6]};
                    end
                    spike_register[i6] = 0;
                    lock6 = 0;
                end
            end
        end

    end
    always @(clear, lock7, spike300, spike301, spike302, spike303, spike304, spike305, spike306, spike307, spike308, spike309, spike310, spike311, spike312, spike313, spike314, spike315, spike316, spike317, spike318, spike319, spike320, spike321, spike322, spike323, spike324, spike325, spike326, spike327, spike328, spike329, spike330, spike331, spike332, spike333, spike334, spike335, spike336, spike337, spike338, spike339, spike340, spike341, spike342, spike343, spike344, spike345, spike346, spike347, spike348, spike349) begin
        spike_register[300] = spike300;

        spike_register[301] = spike301;        spike_register[302] = spike302;        spike_register[303] = spike303;        spike_register[304] = spike304;        spike_register[305] = spike305;        spike_register[306] = spike306;        spike_register[307] = spike307;        spike_register[308] = spike308;        spike_register[309] = spike309;        spike_register[310] = spike310;        spike_register[311] = spike311;        spike_register[312] = spike312;        spike_register[313] = spike313;        spike_register[314] = spike314;        spike_register[315] = spike315;        spike_register[316] = spike316;        spike_register[317] = spike317;        spike_register[318] = spike318;        spike_register[319] = spike319;        spike_register[320] = spike320;        spike_register[321] = spike321;        spike_register[322] = spike322;        spike_register[323] = spike323;        spike_register[324] = spike324;        spike_register[325] = spike325;        spike_register[326] = spike326;        spike_register[327] = spike327;        spike_register[328] = spike328;        spike_register[329] = spike329;        spike_register[330] = spike330;        spike_register[331] = spike331;        spike_register[332] = spike332;        spike_register[333] = spike333;        spike_register[334] = spike334;        spike_register[335] = spike335;        spike_register[336] = spike336;        spike_register[337] = spike337;        spike_register[338] = spike338;        spike_register[339] = spike339;        spike_register[340] = spike340;        spike_register[341] = spike341;        spike_register[342] = spike342;        spike_register[343] = spike343;        spike_register[344] = spike344;        spike_register[345] = spike345;        spike_register[346] = spike346;        spike_register[347] = spike347;        spike_register[348] = spike348;        spike_register[349] = spike349;
        #0.5
        if(clear == 1'b0) begin
            for(i7 = 300; i7 <=349; i7= i7+1) begin
                if(spike_register[i7] == 1 && lock7 == 0) begin
                    lock7 = 1;
                    for(j7 = connection_pointer[i7]; j7 < connection_pointer[i7+1]; j7= j7+1) begin
                        packet7 = #0.1 {neuron_addresses[i7], downstream_connections[j7]};
                    end
                    spike_register[i7] = 0;
                    lock7 = 0;
                end
            end
        end

    end
    always @(clear, lock8, spike350, spike351, spike352, spike353, spike354, spike355, spike356, spike357, spike358, spike359, spike360, spike361, spike362, spike363, spike364, spike365, spike366, spike367, spike368, spike369, spike370, spike371, spike372, spike373, spike374, spike375, spike376, spike377, spike378, spike379, spike380, spike381, spike382, spike383, spike384, spike385, spike386, spike387, spike388, spike389, spike390, spike391, spike392, spike393, spike394, spike395, spike396, spike397, spike398, spike399) begin
        spike_register[350] = spike350;        spike_register[351] = spike351;        spike_register[352] = spike352;        spike_register[353] = spike353;        spike_register[354] = spike354;        spike_register[355] = spike355;        spike_register[356] = spike356;        spike_register[357] = spike357;        spike_register[358] = spike358;        spike_register[359] = spike359;        spike_register[360] = spike360;        spike_register[361] = spike361;        spike_register[362] = spike362;        spike_register[363] = spike363;        spike_register[364] = spike364;        spike_register[365] = spike365;        spike_register[366] = spike366;        spike_register[367] = spike367;        spike_register[368] = spike368;        spike_register[369] = spike369;        spike_register[370] = spike370;        spike_register[371] = spike371;        spike_register[372] = spike372;        spike_register[373] = spike373;        spike_register[374] = spike374;        spike_register[375] = spike375;        spike_register[376] = spike376;        spike_register[377] = spike377;        spike_register[378] = spike378;        spike_register[379] = spike379;        spike_register[380] = spike380;        spike_register[381] = spike381;        spike_register[382] = spike382;        spike_register[383] = spike383;        spike_register[384] = spike384;        spike_register[385] = spike385;        spike_register[386] = spike386;        spike_register[387] = spike387;        spike_register[388] = spike388;        spike_register[389] = spike389;        spike_register[390] = spike390;        spike_register[391] = spike391;        spike_register[392] = spike392;        spike_register[393] = spike393;        spike_register[394] = spike394;        spike_register[395] = spike395;        spike_register[396] = spike396;        spike_register[397] = spike397;        spike_register[398] = spike398;        spike_register[399] = spike399;
        #0.5
        if(clear == 1'b0) begin
            for(i8 = 350; i8 <=399; i8= i8+1) begin
                if(spike_register[i8] == 1 && lock8 == 0) begin
                    lock8 = 1;
                    for(j8 = connection_pointer[i8]; j8 < connection_pointer[i8+1]; j8= j8+1) begin
                        packet8 = #0.1 {neuron_addresses[i8], downstream_connections[j8]};
                    end
                    spike_register[i8] = 0;
                    lock8 = 0;
                end
            end
        end

    end
    always @(clear, lock9, spike400, spike401, spike402, spike403, spike404, spike405, spike406, spike407, spike408, spike409, spike410, spike411, spike412, spike413, spike414, spike415, spike416, spike417, spike418, spike419, spike420, spike421, spike422, spike423, spike424, spike425, spike426, spike427, spike428, spike429, spike430, spike431, spike432, spike433, spike434, spike435, spike436, spike437, spike438, spike439, spike440, spike441, spike442, spike443, spike444, spike445, spike446, spike447, spike448, spike449) begin
        spike_register[400] = spike400;

        spike_register[401] = spike401;        spike_register[402] = spike402;        spike_register[403] = spike403;        spike_register[404] = spike404;        spike_register[405] = spike405;        spike_register[406] = spike406;        spike_register[407] = spike407;        spike_register[408] = spike408;        spike_register[409] = spike409;        spike_register[410] = spike410;        spike_register[411] = spike411;        spike_register[412] = spike412;        spike_register[413] = spike413;        spike_register[414] = spike414;        spike_register[415] = spike415;        spike_register[416] = spike416;        spike_register[417] = spike417;        spike_register[418] = spike418;        spike_register[419] = spike419;        spike_register[420] = spike420;        spike_register[421] = spike421;        spike_register[422] = spike422;        spike_register[423] = spike423;        spike_register[424] = spike424;        spike_register[425] = spike425;        spike_register[426] = spike426;        spike_register[427] = spike427;        spike_register[428] = spike428;        spike_register[429] = spike429;        spike_register[430] = spike430;        spike_register[431] = spike431;        spike_register[432] = spike432;        spike_register[433] = spike433;        spike_register[434] = spike434;        spike_register[435] = spike435;        spike_register[436] = spike436;        spike_register[437] = spike437;        spike_register[438] = spike438;        spike_register[439] = spike439;        spike_register[440] = spike440;        spike_register[441] = spike441;        spike_register[442] = spike442;        spike_register[443] = spike443;        spike_register[444] = spike444;        spike_register[445] = spike445;        spike_register[446] = spike446;        spike_register[447] = spike447;        spike_register[448] = spike448;        spike_register[449] = spike449;
        #0.5
        if(clear == 1'b0) begin
            for(i9 = 400; i9 <=449; i9= i9+1) begin
                if(spike_register[i9] == 1 && lock9 == 0) begin
                    lock9 = 1;
                    for(j9 = connection_pointer[i9]; j9 < connection_pointer[i9+1]; j9= j9+1) begin
                        packet9 = #0.1 {neuron_addresses[i9], downstream_connections[j9]};
                    end
                    spike_register[i9] = 0;
                    lock9 = 0;
                end
            end
        end

    end
    always @(clear, lock10, spike450, spike451, spike452, spike453, spike454, spike455, spike456, spike457, spike458, spike459, spike460, spike461, spike462, spike463, spike464, spike465, spike466, spike467, spike468, spike469, spike470, spike471, spike472, spike473, spike474, spike475, spike476, spike477, spike478, spike479, spike480, spike481, spike482, spike483, spike484, spike485, spike486, spike487, spike488, spike489, spike490, spike491, spike492, spike493, spike494, spike495, spike496, spike497, spike498, spike499) begin
        spike_register[450] = spike450;        spike_register[451] = spike451;        spike_register[452] = spike452;        spike_register[453] = spike453;        spike_register[454] = spike454;        spike_register[455] = spike455;        spike_register[456] = spike456;        spike_register[457] = spike457;        spike_register[458] = spike458;        spike_register[459] = spike459;        spike_register[460] = spike460;        spike_register[461] = spike461;        spike_register[462] = spike462;        spike_register[463] = spike463;        spike_register[464] = spike464;        spike_register[465] = spike465;        spike_register[466] = spike466;        spike_register[467] = spike467;        spike_register[468] = spike468;        spike_register[469] = spike469;        spike_register[470] = spike470;        spike_register[471] = spike471;        spike_register[472] = spike472;        spike_register[473] = spike473;        spike_register[474] = spike474;        spike_register[475] = spike475;        spike_register[476] = spike476;        spike_register[477] = spike477;        spike_register[478] = spike478;        spike_register[479] = spike479;        spike_register[480] = spike480;        spike_register[481] = spike481;        spike_register[482] = spike482;        spike_register[483] = spike483;        spike_register[484] = spike484;        spike_register[485] = spike485;        spike_register[486] = spike486;        spike_register[487] = spike487;        spike_register[488] = spike488;        spike_register[489] = spike489;        spike_register[490] = spike490;        spike_register[491] = spike491;        spike_register[492] = spike492;        spike_register[493] = spike493;        spike_register[494] = spike494;        spike_register[495] = spike495;        spike_register[496] = spike496;        spike_register[497] = spike497;        spike_register[498] = spike498;        spike_register[499] = spike499;
        #0.5
        if(clear == 1'b0) begin
            for(i10 = 450; i10 <=499; i10= i10+1) begin
                if(spike_register[i10] == 1 && lock10 == 0) begin
                    lock10 = 1;
                    for(j10 = connection_pointer[i10]; j10 < connection_pointer[i10+1]; j10= j10+1) begin
                        packet10 = #0.1 {neuron_addresses[i10], downstream_connections[j10]};
                    end
                    spike_register[i10] = 0;
                    lock10 = 0;
                end
            end
        end

    end
    always @(clear, lock11, spike500, spike501, spike502, spike503, spike504, spike505, spike506, spike507, spike508, spike509, spike510, spike511, spike512, spike513, spike514, spike515, spike516, spike517, spike518, spike519, spike520, spike521, spike522, spike523, spike524, spike525, spike526, spike527, spike528, spike529, spike530, spike531, spike532, spike533, spike534, spike535, spike536, spike537, spike538, spike539, spike540, spike541, spike542, spike543, spike544, spike545, spike546, spike547, spike548, spike549) begin
        spike_register[500] = spike500;

        spike_register[501] = spike501;        spike_register[502] = spike502;        spike_register[503] = spike503;        spike_register[504] = spike504;        spike_register[505] = spike505;        spike_register[506] = spike506;        spike_register[507] = spike507;        spike_register[508] = spike508;        spike_register[509] = spike509;        spike_register[510] = spike510;        spike_register[511] = spike511;        spike_register[512] = spike512;        spike_register[513] = spike513;        spike_register[514] = spike514;        spike_register[515] = spike515;        spike_register[516] = spike516;        spike_register[517] = spike517;        spike_register[518] = spike518;        spike_register[519] = spike519;        spike_register[520] = spike520;        spike_register[521] = spike521;        spike_register[522] = spike522;        spike_register[523] = spike523;        spike_register[524] = spike524;        spike_register[525] = spike525;        spike_register[526] = spike526;        spike_register[527] = spike527;        spike_register[528] = spike528;        spike_register[529] = spike529;        spike_register[530] = spike530;        spike_register[531] = spike531;        spike_register[532] = spike532;        spike_register[533] = spike533;        spike_register[534] = spike534;        spike_register[535] = spike535;        spike_register[536] = spike536;        spike_register[537] = spike537;        spike_register[538] = spike538;        spike_register[539] = spike539;        spike_register[540] = spike540;        spike_register[541] = spike541;        spike_register[542] = spike542;        spike_register[543] = spike543;        spike_register[544] = spike544;        spike_register[545] = spike545;        spike_register[546] = spike546;        spike_register[547] = spike547;        spike_register[548] = spike548;        spike_register[549] = spike549;
        #0.5
        if(clear == 1'b0) begin
            for(i11 = 500; i11 <=549; i11= i11+1) begin
                if(spike_register[i11] == 1 && lock11 == 0) begin
                    lock11 = 1;
                    for(j11 = connection_pointer[i11]; j11 < connection_pointer[i11+1]; j11= j11+1) begin
                        packet11 = #0.1 {neuron_addresses[i11], downstream_connections[j11]};
                    end
                    spike_register[i11] = 0;
                    lock11 = 0;
                end
            end
        end

    end
    always @(clear, lock12, spike550, spike551, spike552, spike553, spike554, spike555, spike556, spike557, spike558, spike559, spike560, spike561, spike562, spike563, spike564, spike565, spike566, spike567, spike568, spike569, spike570, spike571, spike572, spike573, spike574, spike575, spike576, spike577, spike578, spike579, spike580, spike581, spike582, spike583, spike584, spike585, spike586, spike587, spike588, spike589, spike590, spike591, spike592, spike593, spike594, spike595, spike596, spike597, spike598, spike599) begin
        spike_register[550] = spike550;        spike_register[551] = spike551;        spike_register[552] = spike552;        spike_register[553] = spike553;        spike_register[554] = spike554;        spike_register[555] = spike555;        spike_register[556] = spike556;        spike_register[557] = spike557;        spike_register[558] = spike558;        spike_register[559] = spike559;        spike_register[560] = spike560;        spike_register[561] = spike561;        spike_register[562] = spike562;        spike_register[563] = spike563;        spike_register[564] = spike564;        spike_register[565] = spike565;        spike_register[566] = spike566;        spike_register[567] = spike567;        spike_register[568] = spike568;        spike_register[569] = spike569;        spike_register[570] = spike570;        spike_register[571] = spike571;        spike_register[572] = spike572;        spike_register[573] = spike573;        spike_register[574] = spike574;        spike_register[575] = spike575;        spike_register[576] = spike576;        spike_register[577] = spike577;        spike_register[578] = spike578;        spike_register[579] = spike579;        spike_register[580] = spike580;        spike_register[581] = spike581;        spike_register[582] = spike582;        spike_register[583] = spike583;        spike_register[584] = spike584;        spike_register[585] = spike585;        spike_register[586] = spike586;        spike_register[587] = spike587;        spike_register[588] = spike588;        spike_register[589] = spike589;        spike_register[590] = spike590;        spike_register[591] = spike591;        spike_register[592] = spike592;        spike_register[593] = spike593;        spike_register[594] = spike594;        spike_register[595] = spike595;        spike_register[596] = spike596;        spike_register[597] = spike597;        spike_register[598] = spike598;        spike_register[599] = spike599;
        #0.5
        if(clear == 1'b0) begin
            for(i12 = 550; i12 <=599; i12= i12+1) begin
                if(spike_register[i12] == 1 && lock12 == 0) begin
                    lock12 = 1;
                    for(j12 = connection_pointer[i12]; j12 < connection_pointer[i12+1]; j12= j12+1) begin
                        packet12 = #0.1 {neuron_addresses[i12], downstream_connections[j12]};
                    end
                    spike_register[i12] = 0;
                    lock12 = 0;
                end
            end
        end

    end
    always @(clear, lock13, spike600, spike601, spike602, spike603, spike604, spike605, spike606, spike607, spike608, spike609, spike610, spike611, spike612, spike613, spike614, spike615, spike616, spike617, spike618, spike619, spike620, spike621, spike622, spike623, spike624, spike625, spike626, spike627, spike628, spike629, spike630, spike631, spike632, spike633, spike634, spike635, spike636, spike637, spike638, spike639, spike640, spike641, spike642, spike643, spike644, spike645, spike646, spike647, spike648, spike649) begin
        spike_register[600] = spike600;

        spike_register[601] = spike601;        spike_register[602] = spike602;        spike_register[603] = spike603;        spike_register[604] = spike604;        spike_register[605] = spike605;        spike_register[606] = spike606;        spike_register[607] = spike607;        spike_register[608] = spike608;        spike_register[609] = spike609;        spike_register[610] = spike610;        spike_register[611] = spike611;        spike_register[612] = spike612;        spike_register[613] = spike613;        spike_register[614] = spike614;        spike_register[615] = spike615;        spike_register[616] = spike616;        spike_register[617] = spike617;        spike_register[618] = spike618;        spike_register[619] = spike619;        spike_register[620] = spike620;        spike_register[621] = spike621;        spike_register[622] = spike622;        spike_register[623] = spike623;        spike_register[624] = spike624;        spike_register[625] = spike625;        spike_register[626] = spike626;        spike_register[627] = spike627;        spike_register[628] = spike628;        spike_register[629] = spike629;        spike_register[630] = spike630;        spike_register[631] = spike631;        spike_register[632] = spike632;        spike_register[633] = spike633;        spike_register[634] = spike634;        spike_register[635] = spike635;        spike_register[636] = spike636;        spike_register[637] = spike637;        spike_register[638] = spike638;        spike_register[639] = spike639;        spike_register[640] = spike640;        spike_register[641] = spike641;        spike_register[642] = spike642;        spike_register[643] = spike643;        spike_register[644] = spike644;        spike_register[645] = spike645;        spike_register[646] = spike646;        spike_register[647] = spike647;        spike_register[648] = spike648;        spike_register[649] = spike649;
        #0.5
        if(clear == 1'b0) begin
            for(i13 = 600; i13 <=649; i13= i13+1) begin
                if(spike_register[i13] == 1 && lock13 == 0) begin
                    lock13 = 1;
                    for(j13 = connection_pointer[i13]; j13 < connection_pointer[i13+1]; j13= j13+1) begin
                        packet13 = #0.1 {neuron_addresses[i13], downstream_connections[j13]};
                    end
                    spike_register[i13] = 0;
                    lock13 = 0;
                end
            end
        end

    end
    always @(clear, lock14, spike650, spike651, spike652, spike653, spike654, spike655, spike656, spike657, spike658, spike659, spike660, spike661, spike662, spike663, spike664, spike665, spike666, spike667, spike668, spike669, spike670, spike671, spike672, spike673, spike674, spike675, spike676, spike677, spike678, spike679, spike680, spike681, spike682, spike683, spike684, spike685, spike686, spike687, spike688, spike689, spike690, spike691, spike692, spike693, spike694, spike695, spike696, spike697, spike698, spike699) begin
        spike_register[650] = spike650;        spike_register[651] = spike651;        spike_register[652] = spike652;        spike_register[653] = spike653;        spike_register[654] = spike654;        spike_register[655] = spike655;        spike_register[656] = spike656;        spike_register[657] = spike657;        spike_register[658] = spike658;        spike_register[659] = spike659;        spike_register[660] = spike660;        spike_register[661] = spike661;        spike_register[662] = spike662;        spike_register[663] = spike663;        spike_register[664] = spike664;        spike_register[665] = spike665;        spike_register[666] = spike666;        spike_register[667] = spike667;        spike_register[668] = spike668;        spike_register[669] = spike669;        spike_register[670] = spike670;        spike_register[671] = spike671;        spike_register[672] = spike672;        spike_register[673] = spike673;        spike_register[674] = spike674;        spike_register[675] = spike675;        spike_register[676] = spike676;        spike_register[677] = spike677;        spike_register[678] = spike678;        spike_register[679] = spike679;        spike_register[680] = spike680;        spike_register[681] = spike681;        spike_register[682] = spike682;        spike_register[683] = spike683;        spike_register[684] = spike684;        spike_register[685] = spike685;        spike_register[686] = spike686;        spike_register[687] = spike687;        spike_register[688] = spike688;        spike_register[689] = spike689;        spike_register[690] = spike690;        spike_register[691] = spike691;        spike_register[692] = spike692;        spike_register[693] = spike693;        spike_register[694] = spike694;        spike_register[695] = spike695;        spike_register[696] = spike696;        spike_register[697] = spike697;        spike_register[698] = spike698;        spike_register[699] = spike699;
        #0.5
        if(clear == 1'b0) begin
            for(i14 = 650; i14 <=699; i14= i14+1) begin
                if(spike_register[i14] == 1 && lock14 == 0) begin
                    lock14 = 1;
                    for(j14 = connection_pointer[i14]; j14 < connection_pointer[i14+1]; j14= j14+1) begin
                        packet14 = #0.1 {neuron_addresses[i14], downstream_connections[j14]};
                    end
                    spike_register[i14] = 0;
                    lock14 = 0;
                end
            end
        end

    end
    always @(clear, lock15, spike700, spike701, spike702, spike703, spike704, spike705, spike706, spike707, spike708, spike709, spike710, spike711, spike712, spike713, spike714, spike715, spike716, spike717, spike718, spike719, spike720, spike721, spike722, spike723, spike724, spike725, spike726, spike727, spike728, spike729, spike730, spike731, spike732, spike733, spike734, spike735, spike736, spike737, spike738, spike739, spike740, spike741, spike742, spike743, spike744, spike745, spike746, spike747, spike748, spike749) begin
        spike_register[700] = spike700;

        spike_register[701] = spike701;        spike_register[702] = spike702;        spike_register[703] = spike703;        spike_register[704] = spike704;        spike_register[705] = spike705;        spike_register[706] = spike706;        spike_register[707] = spike707;        spike_register[708] = spike708;        spike_register[709] = spike709;        spike_register[710] = spike710;        spike_register[711] = spike711;        spike_register[712] = spike712;        spike_register[713] = spike713;        spike_register[714] = spike714;        spike_register[715] = spike715;        spike_register[716] = spike716;        spike_register[717] = spike717;        spike_register[718] = spike718;        spike_register[719] = spike719;        spike_register[720] = spike720;        spike_register[721] = spike721;        spike_register[722] = spike722;        spike_register[723] = spike723;        spike_register[724] = spike724;        spike_register[725] = spike725;        spike_register[726] = spike726;        spike_register[727] = spike727;        spike_register[728] = spike728;        spike_register[729] = spike729;        spike_register[730] = spike730;        spike_register[731] = spike731;        spike_register[732] = spike732;        spike_register[733] = spike733;        spike_register[734] = spike734;        spike_register[735] = spike735;        spike_register[736] = spike736;        spike_register[737] = spike737;        spike_register[738] = spike738;        spike_register[739] = spike739;        spike_register[740] = spike740;        spike_register[741] = spike741;        spike_register[742] = spike742;        spike_register[743] = spike743;        spike_register[744] = spike744;        spike_register[745] = spike745;        spike_register[746] = spike746;        spike_register[747] = spike747;        spike_register[748] = spike748;        spike_register[749] = spike749;
        #0.5
        if(clear == 1'b0) begin
            for(i15 = 700; i15 <=749; i15= i15+1) begin
                if(spike_register[i15] == 1 && lock15 == 0) begin
                    lock15 = 1;
                    for(j15 = connection_pointer[i15]; j15 < connection_pointer[i15+1]; j15= j15+1) begin
                        packet15 = #0.1 {neuron_addresses[i15], downstream_connections[j15]};
                    end
                    spike_register[i15] = 0;
                    lock15 = 0;
                end
            end
        end

    end
    always @(clear, lock16, spike750, spike751, spike752, spike753, spike754, spike755, spike756, spike757, spike758, spike759, spike760, spike761, spike762, spike763, spike764, spike765, spike766, spike767, spike768, spike769, spike770, spike771, spike772, spike773, spike774, spike775, spike776, spike777, spike778, spike779, spike780, spike781, spike782, spike783, spike784, spike785, spike786, spike787, spike788, spike789, spike790, spike791, spike792, spike793, spike794, spike795, spike796, spike797, spike798, spike799) begin
        spike_register[750] = spike750;        spike_register[751] = spike751;        spike_register[752] = spike752;        spike_register[753] = spike753;        spike_register[754] = spike754;        spike_register[755] = spike755;        spike_register[756] = spike756;        spike_register[757] = spike757;        spike_register[758] = spike758;        spike_register[759] = spike759;        spike_register[760] = spike760;        spike_register[761] = spike761;        spike_register[762] = spike762;        spike_register[763] = spike763;        spike_register[764] = spike764;        spike_register[765] = spike765;        spike_register[766] = spike766;        spike_register[767] = spike767;        spike_register[768] = spike768;        spike_register[769] = spike769;        spike_register[770] = spike770;        spike_register[771] = spike771;        spike_register[772] = spike772;        spike_register[773] = spike773;        spike_register[774] = spike774;        spike_register[775] = spike775;        spike_register[776] = spike776;        spike_register[777] = spike777;        spike_register[778] = spike778;        spike_register[779] = spike779;        spike_register[780] = spike780;        spike_register[781] = spike781;        spike_register[782] = spike782;        spike_register[783] = spike783;        spike_register[784] = spike784;        spike_register[785] = spike785;        spike_register[786] = spike786;        spike_register[787] = spike787;        spike_register[788] = spike788;        spike_register[789] = spike789;        spike_register[790] = spike790;        spike_register[791] = spike791;        spike_register[792] = spike792;        spike_register[793] = spike793;        spike_register[794] = spike794;        spike_register[795] = spike795;        spike_register[796] = spike796;        spike_register[797] = spike797;        spike_register[798] = spike798;        spike_register[799] = spike799;
        #0.5
        if(clear == 1'b0) begin
            for(i16 = 750; i16 <=799; i16= i16+1) begin
                if(spike_register[i16] == 1 && lock16 == 0) begin
                    lock16 = 1;
                    for(j16 = connection_pointer[i16]; j16 < connection_pointer[i16+1]; j16= j16+1) begin
                        packet16 = #0.1 {neuron_addresses[i16], downstream_connections[j16]};
                    end
                    spike_register[i16] = 0;
                    lock16 = 0;
                end
            end
        end

    end
    always @(clear, lock17, spike800, spike801, spike802, spike803, spike804, spike805, spike806, spike807, spike808, spike809, spike810, spike811, spike812, spike813, spike814, spike815, spike816, spike817, spike818, spike819, spike820, spike821, spike822, spike823, spike824, spike825, spike826, spike827, spike828, spike829, spike830, spike831, spike832, spike833, spike834, spike835, spike836, spike837, spike838, spike839, spike840, spike841, spike842, spike843, spike844, spike845, spike846, spike847, spike848, spike849) begin
        spike_register[800] = spike800;

        spike_register[801] = spike801;        spike_register[802] = spike802;        spike_register[803] = spike803;        spike_register[804] = spike804;        spike_register[805] = spike805;        spike_register[806] = spike806;        spike_register[807] = spike807;        spike_register[808] = spike808;        spike_register[809] = spike809;        spike_register[810] = spike810;        spike_register[811] = spike811;        spike_register[812] = spike812;        spike_register[813] = spike813;        spike_register[814] = spike814;        spike_register[815] = spike815;        spike_register[816] = spike816;        spike_register[817] = spike817;        spike_register[818] = spike818;        spike_register[819] = spike819;        spike_register[820] = spike820;        spike_register[821] = spike821;        spike_register[822] = spike822;        spike_register[823] = spike823;        spike_register[824] = spike824;        spike_register[825] = spike825;        spike_register[826] = spike826;        spike_register[827] = spike827;        spike_register[828] = spike828;        spike_register[829] = spike829;        spike_register[830] = spike830;        spike_register[831] = spike831;        spike_register[832] = spike832;        spike_register[833] = spike833;        spike_register[834] = spike834;        spike_register[835] = spike835;        spike_register[836] = spike836;        spike_register[837] = spike837;        spike_register[838] = spike838;        spike_register[839] = spike839;        spike_register[840] = spike840;        spike_register[841] = spike841;        spike_register[842] = spike842;        spike_register[843] = spike843;        spike_register[844] = spike844;        spike_register[845] = spike845;        spike_register[846] = spike846;        spike_register[847] = spike847;        spike_register[848] = spike848;        spike_register[849] = spike849;
        #0.5
        if(clear == 1'b0) begin
            for(i17 = 800; i17 <=849; i17= i17+1) begin
                if(spike_register[i17] == 1 && lock17 == 0) begin
                    lock17 = 1;
                    for(j17 = connection_pointer[i17]; j17 < connection_pointer[i17+1]; j17= j17+1) begin
                        packet17 = #0.1 {neuron_addresses[i17], downstream_connections[j17]};
                    end
                    spike_register[i17] = 0;
                    lock17 = 0;
                end
            end
        end

    end
    always @(clear, lock18, spike850, spike851, spike852, spike853, spike854, spike855, spike856, spike857, spike858, spike859, spike860, spike861, spike862, spike863, spike864, spike865, spike866, spike867, spike868, spike869, spike870, spike871, spike872, spike873, spike874, spike875, spike876, spike877, spike878, spike879, spike880, spike881, spike882, spike883, spike884, spike885, spike886, spike887, spike888, spike889, spike890, spike891, spike892, spike893, spike894, spike895, spike896, spike897, spike898, spike899) begin
        spike_register[850] = spike850;        spike_register[851] = spike851;        spike_register[852] = spike852;        spike_register[853] = spike853;        spike_register[854] = spike854;        spike_register[855] = spike855;        spike_register[856] = spike856;        spike_register[857] = spike857;        spike_register[858] = spike858;        spike_register[859] = spike859;        spike_register[860] = spike860;        spike_register[861] = spike861;        spike_register[862] = spike862;        spike_register[863] = spike863;        spike_register[864] = spike864;        spike_register[865] = spike865;        spike_register[866] = spike866;        spike_register[867] = spike867;        spike_register[868] = spike868;        spike_register[869] = spike869;        spike_register[870] = spike870;        spike_register[871] = spike871;        spike_register[872] = spike872;        spike_register[873] = spike873;        spike_register[874] = spike874;        spike_register[875] = spike875;        spike_register[876] = spike876;        spike_register[877] = spike877;        spike_register[878] = spike878;        spike_register[879] = spike879;        spike_register[880] = spike880;        spike_register[881] = spike881;        spike_register[882] = spike882;        spike_register[883] = spike883;        spike_register[884] = spike884;        spike_register[885] = spike885;        spike_register[886] = spike886;        spike_register[887] = spike887;        spike_register[888] = spike888;        spike_register[889] = spike889;        spike_register[890] = spike890;        spike_register[891] = spike891;        spike_register[892] = spike892;        spike_register[893] = spike893;        spike_register[894] = spike894;        spike_register[895] = spike895;        spike_register[896] = spike896;        spike_register[897] = spike897;        spike_register[898] = spike898;        spike_register[899] = spike899;
        #0.5
        if(clear == 1'b0) begin
            for(i18 = 850; i18 <=899; i18= i18+1) begin
                if(spike_register[i18] == 1 && lock18 == 0) begin
                    lock18 = 1;
                    for(j18 = connection_pointer[i18]; j18 < connection_pointer[i18+1]; j18= j18+1) begin
                        packet18 = #0.1 {neuron_addresses[i18], downstream_connections[j18]};
                    end
                    spike_register[i18] = 0;
                    lock18 = 0;
                end
            end
        end

    end
    always @(clear, lock19, spike900, spike901, spike902, spike903, spike904, spike905, spike906, spike907, spike908, spike909, spike910, spike911, spike912, spike913, spike914, spike915, spike916, spike917, spike918, spike919, spike920, spike921, spike922, spike923, spike924, spike925, spike926, spike927, spike928, spike929, spike930, spike931, spike932, spike933, spike934, spike935, spike936, spike937, spike938, spike939, spike940, spike941, spike942, spike943, spike944, spike945, spike946, spike947, spike948, spike949) begin
        spike_register[900] = spike900;

        spike_register[901] = spike901;        spike_register[902] = spike902;        spike_register[903] = spike903;        spike_register[904] = spike904;        spike_register[905] = spike905;        spike_register[906] = spike906;        spike_register[907] = spike907;        spike_register[908] = spike908;        spike_register[909] = spike909;        spike_register[910] = spike910;        spike_register[911] = spike911;        spike_register[912] = spike912;        spike_register[913] = spike913;        spike_register[914] = spike914;        spike_register[915] = spike915;        spike_register[916] = spike916;        spike_register[917] = spike917;        spike_register[918] = spike918;        spike_register[919] = spike919;        spike_register[920] = spike920;        spike_register[921] = spike921;        spike_register[922] = spike922;        spike_register[923] = spike923;        spike_register[924] = spike924;        spike_register[925] = spike925;        spike_register[926] = spike926;        spike_register[927] = spike927;        spike_register[928] = spike928;        spike_register[929] = spike929;        spike_register[930] = spike930;        spike_register[931] = spike931;        spike_register[932] = spike932;        spike_register[933] = spike933;        spike_register[934] = spike934;        spike_register[935] = spike935;        spike_register[936] = spike936;        spike_register[937] = spike937;        spike_register[938] = spike938;        spike_register[939] = spike939;        spike_register[940] = spike940;        spike_register[941] = spike941;        spike_register[942] = spike942;        spike_register[943] = spike943;        spike_register[944] = spike944;        spike_register[945] = spike945;        spike_register[946] = spike946;        spike_register[947] = spike947;        spike_register[948] = spike948;        spike_register[949] = spike949;
        #0.5
        if(clear == 1'b0) begin
            for(i19 = 900; i19 <=949; i19= i19+1) begin
                if(spike_register[i19] == 1 && lock19 == 0) begin
                    lock19 = 1;
                    for(j19 = connection_pointer[i19]; j19 < connection_pointer[i19+1]; j19= j19+1) begin
                        packet19 = #0.1 {neuron_addresses[i19], downstream_connections[j19]};
                    end
                    spike_register[i19] = 0;
                    lock19 = 0;
                end
            end
        end

    end
    always @(clear, lock20, spike950, spike951, spike952, spike953, spike954, spike955, spike956, spike957, spike958, spike959, spike960, spike961, spike962, spike963, spike964, spike965, spike966, spike967, spike968, spike969, spike970, spike971, spike972, spike973, spike974, spike975, spike976, spike977, spike978, spike979, spike980, spike981, spike982, spike983, spike984, spike985, spike986, spike987, spike988, spike989, spike990, spike991, spike992, spike993, spike994, spike995, spike996, spike997, spike998, spike999) begin
        spike_register[950] = spike950;        spike_register[951] = spike951;        spike_register[952] = spike952;        spike_register[953] = spike953;        spike_register[954] = spike954;        spike_register[955] = spike955;        spike_register[956] = spike956;        spike_register[957] = spike957;        spike_register[958] = spike958;        spike_register[959] = spike959;        spike_register[960] = spike960;        spike_register[961] = spike961;        spike_register[962] = spike962;        spike_register[963] = spike963;        spike_register[964] = spike964;        spike_register[965] = spike965;        spike_register[966] = spike966;        spike_register[967] = spike967;        spike_register[968] = spike968;        spike_register[969] = spike969;        spike_register[970] = spike970;        spike_register[971] = spike971;        spike_register[972] = spike972;        spike_register[973] = spike973;        spike_register[974] = spike974;        spike_register[975] = spike975;        spike_register[976] = spike976;        spike_register[977] = spike977;        spike_register[978] = spike978;        spike_register[979] = spike979;        spike_register[980] = spike980;        spike_register[981] = spike981;        spike_register[982] = spike982;        spike_register[983] = spike983;        spike_register[984] = spike984;        spike_register[985] = spike985;        spike_register[986] = spike986;        spike_register[987] = spike987;        spike_register[988] = spike988;        spike_register[989] = spike989;        spike_register[990] = spike990;        spike_register[991] = spike991;        spike_register[992] = spike992;        spike_register[993] = spike993;        spike_register[994] = spike994;        spike_register[995] = spike995;        spike_register[996] = spike996;        spike_register[997] = spike997;        spike_register[998] = spike998;        spike_register[999] = spike999;
        #0.5
        if(clear == 1'b0) begin
            for(i20 = 950; i20 <=999; i20= i20+1) begin
                if(spike_register[i20] == 1 && lock20 == 0) begin
                    lock20 = 1;
                    for(j20 = connection_pointer[i20]; j20 < connection_pointer[i20+1]; j20= j20+1) begin
                        packet20 = #0.1 {neuron_addresses[i20], downstream_connections[j20]};
                    end
                    spike_register[i20] = 0;
                    lock20 = 0;
                end
            end
        end

    end
    always @(clear, lock21, spike1000, spike1001, spike1002, spike1003, spike1004, spike1005, spike1006, spike1007, spike1008, spike1009, spike1010, spike1011, spike1012, spike1013, spike1014, spike1015, spike1016, spike1017, spike1018, spike1019, spike1020, spike1021, spike1022, spike1023) begin
        spike_register[1000] = spike1000;

        spike_register[1001] = spike1001;        spike_register[1002] = spike1002;        spike_register[1003] = spike1003;        spike_register[1004] = spike1004;        spike_register[1005] = spike1005;        spike_register[1006] = spike1006;        spike_register[1007] = spike1007;        spike_register[1008] = spike1008;        spike_register[1009] = spike1009;        spike_register[1010] = spike1010;        spike_register[1011] = spike1011;        spike_register[1012] = spike1012;        spike_register[1013] = spike1013;        spike_register[1014] = spike1014;        spike_register[1015] = spike1015;        spike_register[1016] = spike1016;        spike_register[1017] = spike1017;        spike_register[1018] = spike1018;        spike_register[1019] = spike1019;        spike_register[1020] = spike1020;        spike_register[1021] = spike1021;        spike_register[1022] = spike1022;        spike_register[1023] = spike1023;
        #0.5
        if(clear == 1'b0) begin
            for(i21 = 1000; i21 <=1049; i21= i21+1) begin
                if(spike_register[i21] == 1 && lock21 == 0) begin
                    lock21 = 1;
                    for(j21 = connection_pointer[i21]; j21 < connection_pointer[i21+1]; j21= j21+1) begin
                        packet21 = #0.1 {neuron_addresses[i21], downstream_connections[j21]};
                    end
                    spike_register[i21] = 0;
                    lock21 = 0;
                end
            end
        end

    end
    always @(packet1) begin 
        spike_origin = packet1[23:12];
        spike_destination = packet1[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet2) begin 
        spike_origin = packet2[23:12];
        spike_destination = packet2[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet3) begin 
        spike_origin = packet3[23:12];
        spike_destination = packet3[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet4) begin 
        spike_origin = packet4[23:12];
        spike_destination = packet4[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet5) begin 
        spike_origin = packet5[23:12];
        spike_destination = packet5[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet6) begin 
        spike_origin = packet6[23:12];
        spike_destination = packet6[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet7) begin 
        spike_origin = packet7[23:12];
        spike_destination = packet7[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet8) begin 
        spike_origin = packet8[23:12];
        spike_destination = packet8[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet9) begin 
        spike_origin = packet9[23:12];
        spike_destination = packet9[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet10) begin 
        spike_origin = packet10[23:12];
        spike_destination = packet10[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet11) begin 
        spike_origin = packet11[23:12];
        spike_destination = packet11[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet12) begin 
        spike_origin = packet12[23:12];
        spike_destination = packet12[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet13) begin 
        spike_origin = packet13[23:12];
        spike_destination = packet13[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet14) begin 
        spike_origin = packet14[23:12];
        spike_destination = packet14[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet15) begin 
        spike_origin = packet15[23:12];
        spike_destination = packet15[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet16) begin 
        spike_origin = packet16[23:12];
        spike_destination = packet16[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet17) begin 
        spike_origin = packet17[23:12];
        spike_destination = packet17[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet18) begin 
        spike_origin = packet18[23:12];
        spike_destination = packet18[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet19) begin 
        spike_origin = packet19[23:12];
        spike_destination = packet19[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet20) begin 
        spike_origin = packet20[23:12];
        spike_destination = packet20[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet21) begin 
        spike_origin = packet21[23:12];
        spike_destination = packet21[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(spike_out_source_array[0]) begin 
        spike_out_source0 = spike_out_source_array[0];
    end
    always @(spike_out_source_array[1]) begin 
        spike_out_source1 = spike_out_source_array[1];
    end
    always @(spike_out_source_array[2]) begin 
        spike_out_source2 = spike_out_source_array[2];
    end
    always @(spike_out_source_array[3]) begin 
        spike_out_source3 = spike_out_source_array[3];
    end
    always @(spike_out_source_array[4]) begin 
        spike_out_source4 = spike_out_source_array[4];
    end
    always @(spike_out_source_array[5]) begin 
        spike_out_source5 = spike_out_source_array[5];
    end
    always @(spike_out_source_array[6]) begin 
        spike_out_source6 = spike_out_source_array[6];
    end
    always @(spike_out_source_array[7]) begin 
        spike_out_source7 = spike_out_source_array[7];
    end
    always @(spike_out_source_array[8]) begin 
        spike_out_source8 = spike_out_source_array[8];
    end
    always @(spike_out_source_array[9]) begin 
        spike_out_source9 = spike_out_source_array[9];
    end
    always @(spike_out_source_array[10]) begin 
        spike_out_source10 = spike_out_source_array[10];
    end
    always @(spike_out_source_array[11]) begin 
        spike_out_source11 = spike_out_source_array[11];
    end
    always @(spike_out_source_array[12]) begin 
        spike_out_source12 = spike_out_source_array[12];
    end
    always @(spike_out_source_array[13]) begin 
        spike_out_source13 = spike_out_source_array[13];
    end
    always @(spike_out_source_array[14]) begin 
        spike_out_source14 = spike_out_source_array[14];
    end
    always @(spike_out_source_array[15]) begin 
        spike_out_source15 = spike_out_source_array[15];
    end
    always @(spike_out_source_array[16]) begin 
        spike_out_source16 = spike_out_source_array[16];
    end
    always @(spike_out_source_array[17]) begin 
        spike_out_source17 = spike_out_source_array[17];
    end
    always @(spike_out_source_array[18]) begin 
        spike_out_source18 = spike_out_source_array[18];
    end
    always @(spike_out_source_array[19]) begin 
        spike_out_source19 = spike_out_source_array[19];
    end
    always @(spike_out_source_array[20]) begin 
        spike_out_source20 = spike_out_source_array[20];
    end
    always @(spike_out_source_array[21]) begin 
        spike_out_source21 = spike_out_source_array[21];
    end
    always @(spike_out_source_array[22]) begin 
        spike_out_source22 = spike_out_source_array[22];
    end
    always @(spike_out_source_array[23]) begin 
        spike_out_source23 = spike_out_source_array[23];
    end
    always @(spike_out_source_array[24]) begin 
        spike_out_source24 = spike_out_source_array[24];
    end
    always @(spike_out_source_array[25]) begin 
        spike_out_source25 = spike_out_source_array[25];
    end
    always @(spike_out_source_array[26]) begin 
        spike_out_source26 = spike_out_source_array[26];
    end
    always @(spike_out_source_array[27]) begin 
        spike_out_source27 = spike_out_source_array[27];
    end
    always @(spike_out_source_array[28]) begin 
        spike_out_source28 = spike_out_source_array[28];
    end
    always @(spike_out_source_array[29]) begin 
        spike_out_source29 = spike_out_source_array[29];
    end
    always @(spike_out_source_array[30]) begin 
        spike_out_source30 = spike_out_source_array[30];
    end
    always @(spike_out_source_array[31]) begin 
        spike_out_source31 = spike_out_source_array[31];
    end
    always @(spike_out_source_array[32]) begin 
        spike_out_source32 = spike_out_source_array[32];
    end
    always @(spike_out_source_array[33]) begin 
        spike_out_source33 = spike_out_source_array[33];
    end
    always @(spike_out_source_array[34]) begin 
        spike_out_source34 = spike_out_source_array[34];
    end
    always @(spike_out_source_array[35]) begin 
        spike_out_source35 = spike_out_source_array[35];
    end
    always @(spike_out_source_array[36]) begin 
        spike_out_source36 = spike_out_source_array[36];
    end
    always @(spike_out_source_array[37]) begin 
        spike_out_source37 = spike_out_source_array[37];
    end
    always @(spike_out_source_array[38]) begin 
        spike_out_source38 = spike_out_source_array[38];
    end
    always @(spike_out_source_array[39]) begin 
        spike_out_source39 = spike_out_source_array[39];
    end
    always @(spike_out_source_array[40]) begin 
        spike_out_source40 = spike_out_source_array[40];
    end
    always @(spike_out_source_array[41]) begin 
        spike_out_source41 = spike_out_source_array[41];
    end
    always @(spike_out_source_array[42]) begin 
        spike_out_source42 = spike_out_source_array[42];
    end
    always @(spike_out_source_array[43]) begin 
        spike_out_source43 = spike_out_source_array[43];
    end
    always @(spike_out_source_array[44]) begin 
        spike_out_source44 = spike_out_source_array[44];
    end
    always @(spike_out_source_array[45]) begin 
        spike_out_source45 = spike_out_source_array[45];
    end
    always @(spike_out_source_array[46]) begin 
        spike_out_source46 = spike_out_source_array[46];
    end
    always @(spike_out_source_array[47]) begin 
        spike_out_source47 = spike_out_source_array[47];
    end
    always @(spike_out_source_array[48]) begin 
        spike_out_source48 = spike_out_source_array[48];
    end
    always @(spike_out_source_array[49]) begin 
        spike_out_source49 = spike_out_source_array[49];
    end
    always @(spike_out_source_array[50]) begin 
        spike_out_source50 = spike_out_source_array[50];
    end
    always @(spike_out_source_array[51]) begin 
        spike_out_source51 = spike_out_source_array[51];
    end
    always @(spike_out_source_array[52]) begin 
        spike_out_source52 = spike_out_source_array[52];
    end
    always @(spike_out_source_array[53]) begin 
        spike_out_source53 = spike_out_source_array[53];
    end
    always @(spike_out_source_array[54]) begin 
        spike_out_source54 = spike_out_source_array[54];
    end
    always @(spike_out_source_array[55]) begin 
        spike_out_source55 = spike_out_source_array[55];
    end
    always @(spike_out_source_array[56]) begin 
        spike_out_source56 = spike_out_source_array[56];
    end
    always @(spike_out_source_array[57]) begin 
        spike_out_source57 = spike_out_source_array[57];
    end
    always @(spike_out_source_array[58]) begin 
        spike_out_source58 = spike_out_source_array[58];
    end
    always @(spike_out_source_array[59]) begin 
        spike_out_source59 = spike_out_source_array[59];
    end
    always @(spike_out_source_array[60]) begin 
        spike_out_source60 = spike_out_source_array[60];
    end
    always @(spike_out_source_array[61]) begin 
        spike_out_source61 = spike_out_source_array[61];
    end
    always @(spike_out_source_array[62]) begin 
        spike_out_source62 = spike_out_source_array[62];
    end
    always @(spike_out_source_array[63]) begin 
        spike_out_source63 = spike_out_source_array[63];
    end
    always @(spike_out_source_array[64]) begin 
        spike_out_source64 = spike_out_source_array[64];
    end
    always @(spike_out_source_array[65]) begin 
        spike_out_source65 = spike_out_source_array[65];
    end
    always @(spike_out_source_array[66]) begin 
        spike_out_source66 = spike_out_source_array[66];
    end
    always @(spike_out_source_array[67]) begin 
        spike_out_source67 = spike_out_source_array[67];
    end
    always @(spike_out_source_array[68]) begin 
        spike_out_source68 = spike_out_source_array[68];
    end
    always @(spike_out_source_array[69]) begin 
        spike_out_source69 = spike_out_source_array[69];
    end
    always @(spike_out_source_array[70]) begin 
        spike_out_source70 = spike_out_source_array[70];
    end
    always @(spike_out_source_array[71]) begin 
        spike_out_source71 = spike_out_source_array[71];
    end
    always @(spike_out_source_array[72]) begin 
        spike_out_source72 = spike_out_source_array[72];
    end
    always @(spike_out_source_array[73]) begin 
        spike_out_source73 = spike_out_source_array[73];
    end
    always @(spike_out_source_array[74]) begin 
        spike_out_source74 = spike_out_source_array[74];
    end
    always @(spike_out_source_array[75]) begin 
        spike_out_source75 = spike_out_source_array[75];
    end
    always @(spike_out_source_array[76]) begin 
        spike_out_source76 = spike_out_source_array[76];
    end
    always @(spike_out_source_array[77]) begin 
        spike_out_source77 = spike_out_source_array[77];
    end
    always @(spike_out_source_array[78]) begin 
        spike_out_source78 = spike_out_source_array[78];
    end
    always @(spike_out_source_array[79]) begin 
        spike_out_source79 = spike_out_source_array[79];
    end
    always @(spike_out_source_array[80]) begin 
        spike_out_source80 = spike_out_source_array[80];
    end
    always @(spike_out_source_array[81]) begin 
        spike_out_source81 = spike_out_source_array[81];
    end
    always @(spike_out_source_array[82]) begin 
        spike_out_source82 = spike_out_source_array[82];
    end
    always @(spike_out_source_array[83]) begin 
        spike_out_source83 = spike_out_source_array[83];
    end
    always @(spike_out_source_array[84]) begin 
        spike_out_source84 = spike_out_source_array[84];
    end
    always @(spike_out_source_array[85]) begin 
        spike_out_source85 = spike_out_source_array[85];
    end
    always @(spike_out_source_array[86]) begin 
        spike_out_source86 = spike_out_source_array[86];
    end
    always @(spike_out_source_array[87]) begin 
        spike_out_source87 = spike_out_source_array[87];
    end
    always @(spike_out_source_array[88]) begin 
        spike_out_source88 = spike_out_source_array[88];
    end
    always @(spike_out_source_array[89]) begin 
        spike_out_source89 = spike_out_source_array[89];
    end
    always @(spike_out_source_array[90]) begin 
        spike_out_source90 = spike_out_source_array[90];
    end
    always @(spike_out_source_array[91]) begin 
        spike_out_source91 = spike_out_source_array[91];
    end
    always @(spike_out_source_array[92]) begin 
        spike_out_source92 = spike_out_source_array[92];
    end
    always @(spike_out_source_array[93]) begin 
        spike_out_source93 = spike_out_source_array[93];
    end
    always @(spike_out_source_array[94]) begin 
        spike_out_source94 = spike_out_source_array[94];
    end
    always @(spike_out_source_array[95]) begin 
        spike_out_source95 = spike_out_source_array[95];
    end
    always @(spike_out_source_array[96]) begin 
        spike_out_source96 = spike_out_source_array[96];
    end
    always @(spike_out_source_array[97]) begin 
        spike_out_source97 = spike_out_source_array[97];
    end
    always @(spike_out_source_array[98]) begin 
        spike_out_source98 = spike_out_source_array[98];
    end
    always @(spike_out_source_array[99]) begin 
        spike_out_source99 = spike_out_source_array[99];
    end
    always @(spike_out_source_array[100]) begin 
        spike_out_source100 = spike_out_source_array[100];
    end
    always @(spike_out_source_array[101]) begin 
        spike_out_source101 = spike_out_source_array[101];
    end
    always @(spike_out_source_array[102]) begin 
        spike_out_source102 = spike_out_source_array[102];
    end
    always @(spike_out_source_array[103]) begin 
        spike_out_source103 = spike_out_source_array[103];
    end
    always @(spike_out_source_array[104]) begin 
        spike_out_source104 = spike_out_source_array[104];
    end
    always @(spike_out_source_array[105]) begin 
        spike_out_source105 = spike_out_source_array[105];
    end
    always @(spike_out_source_array[106]) begin 
        spike_out_source106 = spike_out_source_array[106];
    end
    always @(spike_out_source_array[107]) begin 
        spike_out_source107 = spike_out_source_array[107];
    end
    always @(spike_out_source_array[108]) begin 
        spike_out_source108 = spike_out_source_array[108];
    end
    always @(spike_out_source_array[109]) begin 
        spike_out_source109 = spike_out_source_array[109];
    end
    always @(spike_out_source_array[110]) begin 
        spike_out_source110 = spike_out_source_array[110];
    end
    always @(spike_out_source_array[111]) begin 
        spike_out_source111 = spike_out_source_array[111];
    end
    always @(spike_out_source_array[112]) begin 
        spike_out_source112 = spike_out_source_array[112];
    end
    always @(spike_out_source_array[113]) begin 
        spike_out_source113 = spike_out_source_array[113];
    end
    always @(spike_out_source_array[114]) begin 
        spike_out_source114 = spike_out_source_array[114];
    end
    always @(spike_out_source_array[115]) begin 
        spike_out_source115 = spike_out_source_array[115];
    end
    always @(spike_out_source_array[116]) begin 
        spike_out_source116 = spike_out_source_array[116];
    end
    always @(spike_out_source_array[117]) begin 
        spike_out_source117 = spike_out_source_array[117];
    end
    always @(spike_out_source_array[118]) begin 
        spike_out_source118 = spike_out_source_array[118];
    end
    always @(spike_out_source_array[119]) begin 
        spike_out_source119 = spike_out_source_array[119];
    end
    always @(spike_out_source_array[120]) begin 
        spike_out_source120 = spike_out_source_array[120];
    end
    always @(spike_out_source_array[121]) begin 
        spike_out_source121 = spike_out_source_array[121];
    end
    always @(spike_out_source_array[122]) begin 
        spike_out_source122 = spike_out_source_array[122];
    end
    always @(spike_out_source_array[123]) begin 
        spike_out_source123 = spike_out_source_array[123];
    end
    always @(spike_out_source_array[124]) begin 
        spike_out_source124 = spike_out_source_array[124];
    end
    always @(spike_out_source_array[125]) begin 
        spike_out_source125 = spike_out_source_array[125];
    end
    always @(spike_out_source_array[126]) begin 
        spike_out_source126 = spike_out_source_array[126];
    end
    always @(spike_out_source_array[127]) begin 
        spike_out_source127 = spike_out_source_array[127];
    end
    always @(spike_out_source_array[128]) begin 
        spike_out_source128 = spike_out_source_array[128];
    end
    always @(spike_out_source_array[129]) begin 
        spike_out_source129 = spike_out_source_array[129];
    end
    always @(spike_out_source_array[130]) begin 
        spike_out_source130 = spike_out_source_array[130];
    end
    always @(spike_out_source_array[131]) begin 
        spike_out_source131 = spike_out_source_array[131];
    end
    always @(spike_out_source_array[132]) begin 
        spike_out_source132 = spike_out_source_array[132];
    end
    always @(spike_out_source_array[133]) begin 
        spike_out_source133 = spike_out_source_array[133];
    end
    always @(spike_out_source_array[134]) begin 
        spike_out_source134 = spike_out_source_array[134];
    end
    always @(spike_out_source_array[135]) begin 
        spike_out_source135 = spike_out_source_array[135];
    end
    always @(spike_out_source_array[136]) begin 
        spike_out_source136 = spike_out_source_array[136];
    end
    always @(spike_out_source_array[137]) begin 
        spike_out_source137 = spike_out_source_array[137];
    end
    always @(spike_out_source_array[138]) begin 
        spike_out_source138 = spike_out_source_array[138];
    end
    always @(spike_out_source_array[139]) begin 
        spike_out_source139 = spike_out_source_array[139];
    end
    always @(spike_out_source_array[140]) begin 
        spike_out_source140 = spike_out_source_array[140];
    end
    always @(spike_out_source_array[141]) begin 
        spike_out_source141 = spike_out_source_array[141];
    end
    always @(spike_out_source_array[142]) begin 
        spike_out_source142 = spike_out_source_array[142];
    end
    always @(spike_out_source_array[143]) begin 
        spike_out_source143 = spike_out_source_array[143];
    end
    always @(spike_out_source_array[144]) begin 
        spike_out_source144 = spike_out_source_array[144];
    end
    always @(spike_out_source_array[145]) begin 
        spike_out_source145 = spike_out_source_array[145];
    end
    always @(spike_out_source_array[146]) begin 
        spike_out_source146 = spike_out_source_array[146];
    end
    always @(spike_out_source_array[147]) begin 
        spike_out_source147 = spike_out_source_array[147];
    end
    always @(spike_out_source_array[148]) begin 
        spike_out_source148 = spike_out_source_array[148];
    end
    always @(spike_out_source_array[149]) begin 
        spike_out_source149 = spike_out_source_array[149];
    end
    always @(spike_out_source_array[150]) begin 
        spike_out_source150 = spike_out_source_array[150];
    end
    always @(spike_out_source_array[151]) begin 
        spike_out_source151 = spike_out_source_array[151];
    end
    always @(spike_out_source_array[152]) begin 
        spike_out_source152 = spike_out_source_array[152];
    end
    always @(spike_out_source_array[153]) begin 
        spike_out_source153 = spike_out_source_array[153];
    end
    always @(spike_out_source_array[154]) begin 
        spike_out_source154 = spike_out_source_array[154];
    end
    always @(spike_out_source_array[155]) begin 
        spike_out_source155 = spike_out_source_array[155];
    end
    always @(spike_out_source_array[156]) begin 
        spike_out_source156 = spike_out_source_array[156];
    end
    always @(spike_out_source_array[157]) begin 
        spike_out_source157 = spike_out_source_array[157];
    end
    always @(spike_out_source_array[158]) begin 
        spike_out_source158 = spike_out_source_array[158];
    end
    always @(spike_out_source_array[159]) begin 
        spike_out_source159 = spike_out_source_array[159];
    end
    always @(spike_out_source_array[160]) begin 
        spike_out_source160 = spike_out_source_array[160];
    end
    always @(spike_out_source_array[161]) begin 
        spike_out_source161 = spike_out_source_array[161];
    end
    always @(spike_out_source_array[162]) begin 
        spike_out_source162 = spike_out_source_array[162];
    end
    always @(spike_out_source_array[163]) begin 
        spike_out_source163 = spike_out_source_array[163];
    end
    always @(spike_out_source_array[164]) begin 
        spike_out_source164 = spike_out_source_array[164];
    end
    always @(spike_out_source_array[165]) begin 
        spike_out_source165 = spike_out_source_array[165];
    end
    always @(spike_out_source_array[166]) begin 
        spike_out_source166 = spike_out_source_array[166];
    end
    always @(spike_out_source_array[167]) begin 
        spike_out_source167 = spike_out_source_array[167];
    end
    always @(spike_out_source_array[168]) begin 
        spike_out_source168 = spike_out_source_array[168];
    end
    always @(spike_out_source_array[169]) begin 
        spike_out_source169 = spike_out_source_array[169];
    end
    always @(spike_out_source_array[170]) begin 
        spike_out_source170 = spike_out_source_array[170];
    end
    always @(spike_out_source_array[171]) begin 
        spike_out_source171 = spike_out_source_array[171];
    end
    always @(spike_out_source_array[172]) begin 
        spike_out_source172 = spike_out_source_array[172];
    end
    always @(spike_out_source_array[173]) begin 
        spike_out_source173 = spike_out_source_array[173];
    end
    always @(spike_out_source_array[174]) begin 
        spike_out_source174 = spike_out_source_array[174];
    end
    always @(spike_out_source_array[175]) begin 
        spike_out_source175 = spike_out_source_array[175];
    end
    always @(spike_out_source_array[176]) begin 
        spike_out_source176 = spike_out_source_array[176];
    end
    always @(spike_out_source_array[177]) begin 
        spike_out_source177 = spike_out_source_array[177];
    end
    always @(spike_out_source_array[178]) begin 
        spike_out_source178 = spike_out_source_array[178];
    end
    always @(spike_out_source_array[179]) begin 
        spike_out_source179 = spike_out_source_array[179];
    end
    always @(spike_out_source_array[180]) begin 
        spike_out_source180 = spike_out_source_array[180];
    end
    always @(spike_out_source_array[181]) begin 
        spike_out_source181 = spike_out_source_array[181];
    end
    always @(spike_out_source_array[182]) begin 
        spike_out_source182 = spike_out_source_array[182];
    end
    always @(spike_out_source_array[183]) begin 
        spike_out_source183 = spike_out_source_array[183];
    end
    always @(spike_out_source_array[184]) begin 
        spike_out_source184 = spike_out_source_array[184];
    end
    always @(spike_out_source_array[185]) begin 
        spike_out_source185 = spike_out_source_array[185];
    end
    always @(spike_out_source_array[186]) begin 
        spike_out_source186 = spike_out_source_array[186];
    end
    always @(spike_out_source_array[187]) begin 
        spike_out_source187 = spike_out_source_array[187];
    end
    always @(spike_out_source_array[188]) begin 
        spike_out_source188 = spike_out_source_array[188];
    end
    always @(spike_out_source_array[189]) begin 
        spike_out_source189 = spike_out_source_array[189];
    end
    always @(spike_out_source_array[190]) begin 
        spike_out_source190 = spike_out_source_array[190];
    end
    always @(spike_out_source_array[191]) begin 
        spike_out_source191 = spike_out_source_array[191];
    end
    always @(spike_out_source_array[192]) begin 
        spike_out_source192 = spike_out_source_array[192];
    end
    always @(spike_out_source_array[193]) begin 
        spike_out_source193 = spike_out_source_array[193];
    end
    always @(spike_out_source_array[194]) begin 
        spike_out_source194 = spike_out_source_array[194];
    end
    always @(spike_out_source_array[195]) begin 
        spike_out_source195 = spike_out_source_array[195];
    end
    always @(spike_out_source_array[196]) begin 
        spike_out_source196 = spike_out_source_array[196];
    end
    always @(spike_out_source_array[197]) begin 
        spike_out_source197 = spike_out_source_array[197];
    end
    always @(spike_out_source_array[198]) begin 
        spike_out_source198 = spike_out_source_array[198];
    end
    always @(spike_out_source_array[199]) begin 
        spike_out_source199 = spike_out_source_array[199];
    end
    always @(spike_out_source_array[200]) begin 
        spike_out_source200 = spike_out_source_array[200];
    end
    always @(spike_out_source_array[201]) begin 
        spike_out_source201 = spike_out_source_array[201];
    end
    always @(spike_out_source_array[202]) begin 
        spike_out_source202 = spike_out_source_array[202];
    end
    always @(spike_out_source_array[203]) begin 
        spike_out_source203 = spike_out_source_array[203];
    end
    always @(spike_out_source_array[204]) begin 
        spike_out_source204 = spike_out_source_array[204];
    end
    always @(spike_out_source_array[205]) begin 
        spike_out_source205 = spike_out_source_array[205];
    end
    always @(spike_out_source_array[206]) begin 
        spike_out_source206 = spike_out_source_array[206];
    end
    always @(spike_out_source_array[207]) begin 
        spike_out_source207 = spike_out_source_array[207];
    end
    always @(spike_out_source_array[208]) begin 
        spike_out_source208 = spike_out_source_array[208];
    end
    always @(spike_out_source_array[209]) begin 
        spike_out_source209 = spike_out_source_array[209];
    end
    always @(spike_out_source_array[210]) begin 
        spike_out_source210 = spike_out_source_array[210];
    end
    always @(spike_out_source_array[211]) begin 
        spike_out_source211 = spike_out_source_array[211];
    end
    always @(spike_out_source_array[212]) begin 
        spike_out_source212 = spike_out_source_array[212];
    end
    always @(spike_out_source_array[213]) begin 
        spike_out_source213 = spike_out_source_array[213];
    end
    always @(spike_out_source_array[214]) begin 
        spike_out_source214 = spike_out_source_array[214];
    end
    always @(spike_out_source_array[215]) begin 
        spike_out_source215 = spike_out_source_array[215];
    end
    always @(spike_out_source_array[216]) begin 
        spike_out_source216 = spike_out_source_array[216];
    end
    always @(spike_out_source_array[217]) begin 
        spike_out_source217 = spike_out_source_array[217];
    end
    always @(spike_out_source_array[218]) begin 
        spike_out_source218 = spike_out_source_array[218];
    end
    always @(spike_out_source_array[219]) begin 
        spike_out_source219 = spike_out_source_array[219];
    end
    always @(spike_out_source_array[220]) begin 
        spike_out_source220 = spike_out_source_array[220];
    end
    always @(spike_out_source_array[221]) begin 
        spike_out_source221 = spike_out_source_array[221];
    end
    always @(spike_out_source_array[222]) begin 
        spike_out_source222 = spike_out_source_array[222];
    end
    always @(spike_out_source_array[223]) begin 
        spike_out_source223 = spike_out_source_array[223];
    end
    always @(spike_out_source_array[224]) begin 
        spike_out_source224 = spike_out_source_array[224];
    end
    always @(spike_out_source_array[225]) begin 
        spike_out_source225 = spike_out_source_array[225];
    end
    always @(spike_out_source_array[226]) begin 
        spike_out_source226 = spike_out_source_array[226];
    end
    always @(spike_out_source_array[227]) begin 
        spike_out_source227 = spike_out_source_array[227];
    end
    always @(spike_out_source_array[228]) begin 
        spike_out_source228 = spike_out_source_array[228];
    end
    always @(spike_out_source_array[229]) begin 
        spike_out_source229 = spike_out_source_array[229];
    end
    always @(spike_out_source_array[230]) begin 
        spike_out_source230 = spike_out_source_array[230];
    end
    always @(spike_out_source_array[231]) begin 
        spike_out_source231 = spike_out_source_array[231];
    end
    always @(spike_out_source_array[232]) begin 
        spike_out_source232 = spike_out_source_array[232];
    end
    always @(spike_out_source_array[233]) begin 
        spike_out_source233 = spike_out_source_array[233];
    end
    always @(spike_out_source_array[234]) begin 
        spike_out_source234 = spike_out_source_array[234];
    end
    always @(spike_out_source_array[235]) begin 
        spike_out_source235 = spike_out_source_array[235];
    end
    always @(spike_out_source_array[236]) begin 
        spike_out_source236 = spike_out_source_array[236];
    end
    always @(spike_out_source_array[237]) begin 
        spike_out_source237 = spike_out_source_array[237];
    end
    always @(spike_out_source_array[238]) begin 
        spike_out_source238 = spike_out_source_array[238];
    end
    always @(spike_out_source_array[239]) begin 
        spike_out_source239 = spike_out_source_array[239];
    end
    always @(spike_out_source_array[240]) begin 
        spike_out_source240 = spike_out_source_array[240];
    end
    always @(spike_out_source_array[241]) begin 
        spike_out_source241 = spike_out_source_array[241];
    end
    always @(spike_out_source_array[242]) begin 
        spike_out_source242 = spike_out_source_array[242];
    end
    always @(spike_out_source_array[243]) begin 
        spike_out_source243 = spike_out_source_array[243];
    end
    always @(spike_out_source_array[244]) begin 
        spike_out_source244 = spike_out_source_array[244];
    end
    always @(spike_out_source_array[245]) begin 
        spike_out_source245 = spike_out_source_array[245];
    end
    always @(spike_out_source_array[246]) begin 
        spike_out_source246 = spike_out_source_array[246];
    end
    always @(spike_out_source_array[247]) begin 
        spike_out_source247 = spike_out_source_array[247];
    end
    always @(spike_out_source_array[248]) begin 
        spike_out_source248 = spike_out_source_array[248];
    end
    always @(spike_out_source_array[249]) begin 
        spike_out_source249 = spike_out_source_array[249];
    end
    always @(spike_out_source_array[250]) begin 
        spike_out_source250 = spike_out_source_array[250];
    end
    always @(spike_out_source_array[251]) begin 
        spike_out_source251 = spike_out_source_array[251];
    end
    always @(spike_out_source_array[252]) begin 
        spike_out_source252 = spike_out_source_array[252];
    end
    always @(spike_out_source_array[253]) begin 
        spike_out_source253 = spike_out_source_array[253];
    end
    always @(spike_out_source_array[254]) begin 
        spike_out_source254 = spike_out_source_array[254];
    end
    always @(spike_out_source_array[255]) begin 
        spike_out_source255 = spike_out_source_array[255];
    end
    always @(spike_out_source_array[256]) begin 
        spike_out_source256 = spike_out_source_array[256];
    end
    always @(spike_out_source_array[257]) begin 
        spike_out_source257 = spike_out_source_array[257];
    end
    always @(spike_out_source_array[258]) begin 
        spike_out_source258 = spike_out_source_array[258];
    end
    always @(spike_out_source_array[259]) begin 
        spike_out_source259 = spike_out_source_array[259];
    end
    always @(spike_out_source_array[260]) begin 
        spike_out_source260 = spike_out_source_array[260];
    end
    always @(spike_out_source_array[261]) begin 
        spike_out_source261 = spike_out_source_array[261];
    end
    always @(spike_out_source_array[262]) begin 
        spike_out_source262 = spike_out_source_array[262];
    end
    always @(spike_out_source_array[263]) begin 
        spike_out_source263 = spike_out_source_array[263];
    end
    always @(spike_out_source_array[264]) begin 
        spike_out_source264 = spike_out_source_array[264];
    end
    always @(spike_out_source_array[265]) begin 
        spike_out_source265 = spike_out_source_array[265];
    end
    always @(spike_out_source_array[266]) begin 
        spike_out_source266 = spike_out_source_array[266];
    end
    always @(spike_out_source_array[267]) begin 
        spike_out_source267 = spike_out_source_array[267];
    end
    always @(spike_out_source_array[268]) begin 
        spike_out_source268 = spike_out_source_array[268];
    end
    always @(spike_out_source_array[269]) begin 
        spike_out_source269 = spike_out_source_array[269];
    end
    always @(spike_out_source_array[270]) begin 
        spike_out_source270 = spike_out_source_array[270];
    end
    always @(spike_out_source_array[271]) begin 
        spike_out_source271 = spike_out_source_array[271];
    end
    always @(spike_out_source_array[272]) begin 
        spike_out_source272 = spike_out_source_array[272];
    end
    always @(spike_out_source_array[273]) begin 
        spike_out_source273 = spike_out_source_array[273];
    end
    always @(spike_out_source_array[274]) begin 
        spike_out_source274 = spike_out_source_array[274];
    end
    always @(spike_out_source_array[275]) begin 
        spike_out_source275 = spike_out_source_array[275];
    end
    always @(spike_out_source_array[276]) begin 
        spike_out_source276 = spike_out_source_array[276];
    end
    always @(spike_out_source_array[277]) begin 
        spike_out_source277 = spike_out_source_array[277];
    end
    always @(spike_out_source_array[278]) begin 
        spike_out_source278 = spike_out_source_array[278];
    end
    always @(spike_out_source_array[279]) begin 
        spike_out_source279 = spike_out_source_array[279];
    end
    always @(spike_out_source_array[280]) begin 
        spike_out_source280 = spike_out_source_array[280];
    end
    always @(spike_out_source_array[281]) begin 
        spike_out_source281 = spike_out_source_array[281];
    end
    always @(spike_out_source_array[282]) begin 
        spike_out_source282 = spike_out_source_array[282];
    end
    always @(spike_out_source_array[283]) begin 
        spike_out_source283 = spike_out_source_array[283];
    end
    always @(spike_out_source_array[284]) begin 
        spike_out_source284 = spike_out_source_array[284];
    end
    always @(spike_out_source_array[285]) begin 
        spike_out_source285 = spike_out_source_array[285];
    end
    always @(spike_out_source_array[286]) begin 
        spike_out_source286 = spike_out_source_array[286];
    end
    always @(spike_out_source_array[287]) begin 
        spike_out_source287 = spike_out_source_array[287];
    end
    always @(spike_out_source_array[288]) begin 
        spike_out_source288 = spike_out_source_array[288];
    end
    always @(spike_out_source_array[289]) begin 
        spike_out_source289 = spike_out_source_array[289];
    end
    always @(spike_out_source_array[290]) begin 
        spike_out_source290 = spike_out_source_array[290];
    end
    always @(spike_out_source_array[291]) begin 
        spike_out_source291 = spike_out_source_array[291];
    end
    always @(spike_out_source_array[292]) begin 
        spike_out_source292 = spike_out_source_array[292];
    end
    always @(spike_out_source_array[293]) begin 
        spike_out_source293 = spike_out_source_array[293];
    end
    always @(spike_out_source_array[294]) begin 
        spike_out_source294 = spike_out_source_array[294];
    end
    always @(spike_out_source_array[295]) begin 
        spike_out_source295 = spike_out_source_array[295];
    end
    always @(spike_out_source_array[296]) begin 
        spike_out_source296 = spike_out_source_array[296];
    end
    always @(spike_out_source_array[297]) begin 
        spike_out_source297 = spike_out_source_array[297];
    end
    always @(spike_out_source_array[298]) begin 
        spike_out_source298 = spike_out_source_array[298];
    end
    always @(spike_out_source_array[299]) begin 
        spike_out_source299 = spike_out_source_array[299];
    end
    always @(spike_out_source_array[300]) begin 
        spike_out_source300 = spike_out_source_array[300];
    end
    always @(spike_out_source_array[301]) begin 
        spike_out_source301 = spike_out_source_array[301];
    end
    always @(spike_out_source_array[302]) begin 
        spike_out_source302 = spike_out_source_array[302];
    end
    always @(spike_out_source_array[303]) begin 
        spike_out_source303 = spike_out_source_array[303];
    end
    always @(spike_out_source_array[304]) begin 
        spike_out_source304 = spike_out_source_array[304];
    end
    always @(spike_out_source_array[305]) begin 
        spike_out_source305 = spike_out_source_array[305];
    end
    always @(spike_out_source_array[306]) begin 
        spike_out_source306 = spike_out_source_array[306];
    end
    always @(spike_out_source_array[307]) begin 
        spike_out_source307 = spike_out_source_array[307];
    end
    always @(spike_out_source_array[308]) begin 
        spike_out_source308 = spike_out_source_array[308];
    end
    always @(spike_out_source_array[309]) begin 
        spike_out_source309 = spike_out_source_array[309];
    end
    always @(spike_out_source_array[310]) begin 
        spike_out_source310 = spike_out_source_array[310];
    end
    always @(spike_out_source_array[311]) begin 
        spike_out_source311 = spike_out_source_array[311];
    end
    always @(spike_out_source_array[312]) begin 
        spike_out_source312 = spike_out_source_array[312];
    end
    always @(spike_out_source_array[313]) begin 
        spike_out_source313 = spike_out_source_array[313];
    end
    always @(spike_out_source_array[314]) begin 
        spike_out_source314 = spike_out_source_array[314];
    end
    always @(spike_out_source_array[315]) begin 
        spike_out_source315 = spike_out_source_array[315];
    end
    always @(spike_out_source_array[316]) begin 
        spike_out_source316 = spike_out_source_array[316];
    end
    always @(spike_out_source_array[317]) begin 
        spike_out_source317 = spike_out_source_array[317];
    end
    always @(spike_out_source_array[318]) begin 
        spike_out_source318 = spike_out_source_array[318];
    end
    always @(spike_out_source_array[319]) begin 
        spike_out_source319 = spike_out_source_array[319];
    end
    always @(spike_out_source_array[320]) begin 
        spike_out_source320 = spike_out_source_array[320];
    end
    always @(spike_out_source_array[321]) begin 
        spike_out_source321 = spike_out_source_array[321];
    end
    always @(spike_out_source_array[322]) begin 
        spike_out_source322 = spike_out_source_array[322];
    end
    always @(spike_out_source_array[323]) begin 
        spike_out_source323 = spike_out_source_array[323];
    end
    always @(spike_out_source_array[324]) begin 
        spike_out_source324 = spike_out_source_array[324];
    end
    always @(spike_out_source_array[325]) begin 
        spike_out_source325 = spike_out_source_array[325];
    end
    always @(spike_out_source_array[326]) begin 
        spike_out_source326 = spike_out_source_array[326];
    end
    always @(spike_out_source_array[327]) begin 
        spike_out_source327 = spike_out_source_array[327];
    end
    always @(spike_out_source_array[328]) begin 
        spike_out_source328 = spike_out_source_array[328];
    end
    always @(spike_out_source_array[329]) begin 
        spike_out_source329 = spike_out_source_array[329];
    end
    always @(spike_out_source_array[330]) begin 
        spike_out_source330 = spike_out_source_array[330];
    end
    always @(spike_out_source_array[331]) begin 
        spike_out_source331 = spike_out_source_array[331];
    end
    always @(spike_out_source_array[332]) begin 
        spike_out_source332 = spike_out_source_array[332];
    end
    always @(spike_out_source_array[333]) begin 
        spike_out_source333 = spike_out_source_array[333];
    end
    always @(spike_out_source_array[334]) begin 
        spike_out_source334 = spike_out_source_array[334];
    end
    always @(spike_out_source_array[335]) begin 
        spike_out_source335 = spike_out_source_array[335];
    end
    always @(spike_out_source_array[336]) begin 
        spike_out_source336 = spike_out_source_array[336];
    end
    always @(spike_out_source_array[337]) begin 
        spike_out_source337 = spike_out_source_array[337];
    end
    always @(spike_out_source_array[338]) begin 
        spike_out_source338 = spike_out_source_array[338];
    end
    always @(spike_out_source_array[339]) begin 
        spike_out_source339 = spike_out_source_array[339];
    end
    always @(spike_out_source_array[340]) begin 
        spike_out_source340 = spike_out_source_array[340];
    end
    always @(spike_out_source_array[341]) begin 
        spike_out_source341 = spike_out_source_array[341];
    end
    always @(spike_out_source_array[342]) begin 
        spike_out_source342 = spike_out_source_array[342];
    end
    always @(spike_out_source_array[343]) begin 
        spike_out_source343 = spike_out_source_array[343];
    end
    always @(spike_out_source_array[344]) begin 
        spike_out_source344 = spike_out_source_array[344];
    end
    always @(spike_out_source_array[345]) begin 
        spike_out_source345 = spike_out_source_array[345];
    end
    always @(spike_out_source_array[346]) begin 
        spike_out_source346 = spike_out_source_array[346];
    end
    always @(spike_out_source_array[347]) begin 
        spike_out_source347 = spike_out_source_array[347];
    end
    always @(spike_out_source_array[348]) begin 
        spike_out_source348 = spike_out_source_array[348];
    end
    always @(spike_out_source_array[349]) begin 
        spike_out_source349 = spike_out_source_array[349];
    end
    always @(spike_out_source_array[350]) begin 
        spike_out_source350 = spike_out_source_array[350];
    end
    always @(spike_out_source_array[351]) begin 
        spike_out_source351 = spike_out_source_array[351];
    end
    always @(spike_out_source_array[352]) begin 
        spike_out_source352 = spike_out_source_array[352];
    end
    always @(spike_out_source_array[353]) begin 
        spike_out_source353 = spike_out_source_array[353];
    end
    always @(spike_out_source_array[354]) begin 
        spike_out_source354 = spike_out_source_array[354];
    end
    always @(spike_out_source_array[355]) begin 
        spike_out_source355 = spike_out_source_array[355];
    end
    always @(spike_out_source_array[356]) begin 
        spike_out_source356 = spike_out_source_array[356];
    end
    always @(spike_out_source_array[357]) begin 
        spike_out_source357 = spike_out_source_array[357];
    end
    always @(spike_out_source_array[358]) begin 
        spike_out_source358 = spike_out_source_array[358];
    end
    always @(spike_out_source_array[359]) begin 
        spike_out_source359 = spike_out_source_array[359];
    end
    always @(spike_out_source_array[360]) begin 
        spike_out_source360 = spike_out_source_array[360];
    end
    always @(spike_out_source_array[361]) begin 
        spike_out_source361 = spike_out_source_array[361];
    end
    always @(spike_out_source_array[362]) begin 
        spike_out_source362 = spike_out_source_array[362];
    end
    always @(spike_out_source_array[363]) begin 
        spike_out_source363 = spike_out_source_array[363];
    end
    always @(spike_out_source_array[364]) begin 
        spike_out_source364 = spike_out_source_array[364];
    end
    always @(spike_out_source_array[365]) begin 
        spike_out_source365 = spike_out_source_array[365];
    end
    always @(spike_out_source_array[366]) begin 
        spike_out_source366 = spike_out_source_array[366];
    end
    always @(spike_out_source_array[367]) begin 
        spike_out_source367 = spike_out_source_array[367];
    end
    always @(spike_out_source_array[368]) begin 
        spike_out_source368 = spike_out_source_array[368];
    end
    always @(spike_out_source_array[369]) begin 
        spike_out_source369 = spike_out_source_array[369];
    end
    always @(spike_out_source_array[370]) begin 
        spike_out_source370 = spike_out_source_array[370];
    end
    always @(spike_out_source_array[371]) begin 
        spike_out_source371 = spike_out_source_array[371];
    end
    always @(spike_out_source_array[372]) begin 
        spike_out_source372 = spike_out_source_array[372];
    end
    always @(spike_out_source_array[373]) begin 
        spike_out_source373 = spike_out_source_array[373];
    end
    always @(spike_out_source_array[374]) begin 
        spike_out_source374 = spike_out_source_array[374];
    end
    always @(spike_out_source_array[375]) begin 
        spike_out_source375 = spike_out_source_array[375];
    end
    always @(spike_out_source_array[376]) begin 
        spike_out_source376 = spike_out_source_array[376];
    end
    always @(spike_out_source_array[377]) begin 
        spike_out_source377 = spike_out_source_array[377];
    end
    always @(spike_out_source_array[378]) begin 
        spike_out_source378 = spike_out_source_array[378];
    end
    always @(spike_out_source_array[379]) begin 
        spike_out_source379 = spike_out_source_array[379];
    end
    always @(spike_out_source_array[380]) begin 
        spike_out_source380 = spike_out_source_array[380];
    end
    always @(spike_out_source_array[381]) begin 
        spike_out_source381 = spike_out_source_array[381];
    end
    always @(spike_out_source_array[382]) begin 
        spike_out_source382 = spike_out_source_array[382];
    end
    always @(spike_out_source_array[383]) begin 
        spike_out_source383 = spike_out_source_array[383];
    end
    always @(spike_out_source_array[384]) begin 
        spike_out_source384 = spike_out_source_array[384];
    end
    always @(spike_out_source_array[385]) begin 
        spike_out_source385 = spike_out_source_array[385];
    end
    always @(spike_out_source_array[386]) begin 
        spike_out_source386 = spike_out_source_array[386];
    end
    always @(spike_out_source_array[387]) begin 
        spike_out_source387 = spike_out_source_array[387];
    end
    always @(spike_out_source_array[388]) begin 
        spike_out_source388 = spike_out_source_array[388];
    end
    always @(spike_out_source_array[389]) begin 
        spike_out_source389 = spike_out_source_array[389];
    end
    always @(spike_out_source_array[390]) begin 
        spike_out_source390 = spike_out_source_array[390];
    end
    always @(spike_out_source_array[391]) begin 
        spike_out_source391 = spike_out_source_array[391];
    end
    always @(spike_out_source_array[392]) begin 
        spike_out_source392 = spike_out_source_array[392];
    end
    always @(spike_out_source_array[393]) begin 
        spike_out_source393 = spike_out_source_array[393];
    end
    always @(spike_out_source_array[394]) begin 
        spike_out_source394 = spike_out_source_array[394];
    end
    always @(spike_out_source_array[395]) begin 
        spike_out_source395 = spike_out_source_array[395];
    end
    always @(spike_out_source_array[396]) begin 
        spike_out_source396 = spike_out_source_array[396];
    end
    always @(spike_out_source_array[397]) begin 
        spike_out_source397 = spike_out_source_array[397];
    end
    always @(spike_out_source_array[398]) begin 
        spike_out_source398 = spike_out_source_array[398];
    end
    always @(spike_out_source_array[399]) begin 
        spike_out_source399 = spike_out_source_array[399];
    end
    always @(spike_out_source_array[400]) begin 
        spike_out_source400 = spike_out_source_array[400];
    end
    always @(spike_out_source_array[401]) begin 
        spike_out_source401 = spike_out_source_array[401];
    end
    always @(spike_out_source_array[402]) begin 
        spike_out_source402 = spike_out_source_array[402];
    end
    always @(spike_out_source_array[403]) begin 
        spike_out_source403 = spike_out_source_array[403];
    end
    always @(spike_out_source_array[404]) begin 
        spike_out_source404 = spike_out_source_array[404];
    end
    always @(spike_out_source_array[405]) begin 
        spike_out_source405 = spike_out_source_array[405];
    end
    always @(spike_out_source_array[406]) begin 
        spike_out_source406 = spike_out_source_array[406];
    end
    always @(spike_out_source_array[407]) begin 
        spike_out_source407 = spike_out_source_array[407];
    end
    always @(spike_out_source_array[408]) begin 
        spike_out_source408 = spike_out_source_array[408];
    end
    always @(spike_out_source_array[409]) begin 
        spike_out_source409 = spike_out_source_array[409];
    end
    always @(spike_out_source_array[410]) begin 
        spike_out_source410 = spike_out_source_array[410];
    end
    always @(spike_out_source_array[411]) begin 
        spike_out_source411 = spike_out_source_array[411];
    end
    always @(spike_out_source_array[412]) begin 
        spike_out_source412 = spike_out_source_array[412];
    end
    always @(spike_out_source_array[413]) begin 
        spike_out_source413 = spike_out_source_array[413];
    end
    always @(spike_out_source_array[414]) begin 
        spike_out_source414 = spike_out_source_array[414];
    end
    always @(spike_out_source_array[415]) begin 
        spike_out_source415 = spike_out_source_array[415];
    end
    always @(spike_out_source_array[416]) begin 
        spike_out_source416 = spike_out_source_array[416];
    end
    always @(spike_out_source_array[417]) begin 
        spike_out_source417 = spike_out_source_array[417];
    end
    always @(spike_out_source_array[418]) begin 
        spike_out_source418 = spike_out_source_array[418];
    end
    always @(spike_out_source_array[419]) begin 
        spike_out_source419 = spike_out_source_array[419];
    end
    always @(spike_out_source_array[420]) begin 
        spike_out_source420 = spike_out_source_array[420];
    end
    always @(spike_out_source_array[421]) begin 
        spike_out_source421 = spike_out_source_array[421];
    end
    always @(spike_out_source_array[422]) begin 
        spike_out_source422 = spike_out_source_array[422];
    end
    always @(spike_out_source_array[423]) begin 
        spike_out_source423 = spike_out_source_array[423];
    end
    always @(spike_out_source_array[424]) begin 
        spike_out_source424 = spike_out_source_array[424];
    end
    always @(spike_out_source_array[425]) begin 
        spike_out_source425 = spike_out_source_array[425];
    end
    always @(spike_out_source_array[426]) begin 
        spike_out_source426 = spike_out_source_array[426];
    end
    always @(spike_out_source_array[427]) begin 
        spike_out_source427 = spike_out_source_array[427];
    end
    always @(spike_out_source_array[428]) begin 
        spike_out_source428 = spike_out_source_array[428];
    end
    always @(spike_out_source_array[429]) begin 
        spike_out_source429 = spike_out_source_array[429];
    end
    always @(spike_out_source_array[430]) begin 
        spike_out_source430 = spike_out_source_array[430];
    end
    always @(spike_out_source_array[431]) begin 
        spike_out_source431 = spike_out_source_array[431];
    end
    always @(spike_out_source_array[432]) begin 
        spike_out_source432 = spike_out_source_array[432];
    end
    always @(spike_out_source_array[433]) begin 
        spike_out_source433 = spike_out_source_array[433];
    end
    always @(spike_out_source_array[434]) begin 
        spike_out_source434 = spike_out_source_array[434];
    end
    always @(spike_out_source_array[435]) begin 
        spike_out_source435 = spike_out_source_array[435];
    end
    always @(spike_out_source_array[436]) begin 
        spike_out_source436 = spike_out_source_array[436];
    end
    always @(spike_out_source_array[437]) begin 
        spike_out_source437 = spike_out_source_array[437];
    end
    always @(spike_out_source_array[438]) begin 
        spike_out_source438 = spike_out_source_array[438];
    end
    always @(spike_out_source_array[439]) begin 
        spike_out_source439 = spike_out_source_array[439];
    end
    always @(spike_out_source_array[440]) begin 
        spike_out_source440 = spike_out_source_array[440];
    end
    always @(spike_out_source_array[441]) begin 
        spike_out_source441 = spike_out_source_array[441];
    end
    always @(spike_out_source_array[442]) begin 
        spike_out_source442 = spike_out_source_array[442];
    end
    always @(spike_out_source_array[443]) begin 
        spike_out_source443 = spike_out_source_array[443];
    end
    always @(spike_out_source_array[444]) begin 
        spike_out_source444 = spike_out_source_array[444];
    end
    always @(spike_out_source_array[445]) begin 
        spike_out_source445 = spike_out_source_array[445];
    end
    always @(spike_out_source_array[446]) begin 
        spike_out_source446 = spike_out_source_array[446];
    end
    always @(spike_out_source_array[447]) begin 
        spike_out_source447 = spike_out_source_array[447];
    end
    always @(spike_out_source_array[448]) begin 
        spike_out_source448 = spike_out_source_array[448];
    end
    always @(spike_out_source_array[449]) begin 
        spike_out_source449 = spike_out_source_array[449];
    end
    always @(spike_out_source_array[450]) begin 
        spike_out_source450 = spike_out_source_array[450];
    end
    always @(spike_out_source_array[451]) begin 
        spike_out_source451 = spike_out_source_array[451];
    end
    always @(spike_out_source_array[452]) begin 
        spike_out_source452 = spike_out_source_array[452];
    end
    always @(spike_out_source_array[453]) begin 
        spike_out_source453 = spike_out_source_array[453];
    end
    always @(spike_out_source_array[454]) begin 
        spike_out_source454 = spike_out_source_array[454];
    end
    always @(spike_out_source_array[455]) begin 
        spike_out_source455 = spike_out_source_array[455];
    end
    always @(spike_out_source_array[456]) begin 
        spike_out_source456 = spike_out_source_array[456];
    end
    always @(spike_out_source_array[457]) begin 
        spike_out_source457 = spike_out_source_array[457];
    end
    always @(spike_out_source_array[458]) begin 
        spike_out_source458 = spike_out_source_array[458];
    end
    always @(spike_out_source_array[459]) begin 
        spike_out_source459 = spike_out_source_array[459];
    end
    always @(spike_out_source_array[460]) begin 
        spike_out_source460 = spike_out_source_array[460];
    end
    always @(spike_out_source_array[461]) begin 
        spike_out_source461 = spike_out_source_array[461];
    end
    always @(spike_out_source_array[462]) begin 
        spike_out_source462 = spike_out_source_array[462];
    end
    always @(spike_out_source_array[463]) begin 
        spike_out_source463 = spike_out_source_array[463];
    end
    always @(spike_out_source_array[464]) begin 
        spike_out_source464 = spike_out_source_array[464];
    end
    always @(spike_out_source_array[465]) begin 
        spike_out_source465 = spike_out_source_array[465];
    end
    always @(spike_out_source_array[466]) begin 
        spike_out_source466 = spike_out_source_array[466];
    end
    always @(spike_out_source_array[467]) begin 
        spike_out_source467 = spike_out_source_array[467];
    end
    always @(spike_out_source_array[468]) begin 
        spike_out_source468 = spike_out_source_array[468];
    end
    always @(spike_out_source_array[469]) begin 
        spike_out_source469 = spike_out_source_array[469];
    end
    always @(spike_out_source_array[470]) begin 
        spike_out_source470 = spike_out_source_array[470];
    end
    always @(spike_out_source_array[471]) begin 
        spike_out_source471 = spike_out_source_array[471];
    end
    always @(spike_out_source_array[472]) begin 
        spike_out_source472 = spike_out_source_array[472];
    end
    always @(spike_out_source_array[473]) begin 
        spike_out_source473 = spike_out_source_array[473];
    end
    always @(spike_out_source_array[474]) begin 
        spike_out_source474 = spike_out_source_array[474];
    end
    always @(spike_out_source_array[475]) begin 
        spike_out_source475 = spike_out_source_array[475];
    end
    always @(spike_out_source_array[476]) begin 
        spike_out_source476 = spike_out_source_array[476];
    end
    always @(spike_out_source_array[477]) begin 
        spike_out_source477 = spike_out_source_array[477];
    end
    always @(spike_out_source_array[478]) begin 
        spike_out_source478 = spike_out_source_array[478];
    end
    always @(spike_out_source_array[479]) begin 
        spike_out_source479 = spike_out_source_array[479];
    end
    always @(spike_out_source_array[480]) begin 
        spike_out_source480 = spike_out_source_array[480];
    end
    always @(spike_out_source_array[481]) begin 
        spike_out_source481 = spike_out_source_array[481];
    end
    always @(spike_out_source_array[482]) begin 
        spike_out_source482 = spike_out_source_array[482];
    end
    always @(spike_out_source_array[483]) begin 
        spike_out_source483 = spike_out_source_array[483];
    end
    always @(spike_out_source_array[484]) begin 
        spike_out_source484 = spike_out_source_array[484];
    end
    always @(spike_out_source_array[485]) begin 
        spike_out_source485 = spike_out_source_array[485];
    end
    always @(spike_out_source_array[486]) begin 
        spike_out_source486 = spike_out_source_array[486];
    end
    always @(spike_out_source_array[487]) begin 
        spike_out_source487 = spike_out_source_array[487];
    end
    always @(spike_out_source_array[488]) begin 
        spike_out_source488 = spike_out_source_array[488];
    end
    always @(spike_out_source_array[489]) begin 
        spike_out_source489 = spike_out_source_array[489];
    end
    always @(spike_out_source_array[490]) begin 
        spike_out_source490 = spike_out_source_array[490];
    end
    always @(spike_out_source_array[491]) begin 
        spike_out_source491 = spike_out_source_array[491];
    end
    always @(spike_out_source_array[492]) begin 
        spike_out_source492 = spike_out_source_array[492];
    end
    always @(spike_out_source_array[493]) begin 
        spike_out_source493 = spike_out_source_array[493];
    end
    always @(spike_out_source_array[494]) begin 
        spike_out_source494 = spike_out_source_array[494];
    end
    always @(spike_out_source_array[495]) begin 
        spike_out_source495 = spike_out_source_array[495];
    end
    always @(spike_out_source_array[496]) begin 
        spike_out_source496 = spike_out_source_array[496];
    end
    always @(spike_out_source_array[497]) begin 
        spike_out_source497 = spike_out_source_array[497];
    end
    always @(spike_out_source_array[498]) begin 
        spike_out_source498 = spike_out_source_array[498];
    end
    always @(spike_out_source_array[499]) begin 
        spike_out_source499 = spike_out_source_array[499];
    end
    always @(spike_out_source_array[500]) begin 
        spike_out_source500 = spike_out_source_array[500];
    end
    always @(spike_out_source_array[501]) begin 
        spike_out_source501 = spike_out_source_array[501];
    end
    always @(spike_out_source_array[502]) begin 
        spike_out_source502 = spike_out_source_array[502];
    end
    always @(spike_out_source_array[503]) begin 
        spike_out_source503 = spike_out_source_array[503];
    end
    always @(spike_out_source_array[504]) begin 
        spike_out_source504 = spike_out_source_array[504];
    end
    always @(spike_out_source_array[505]) begin 
        spike_out_source505 = spike_out_source_array[505];
    end
    always @(spike_out_source_array[506]) begin 
        spike_out_source506 = spike_out_source_array[506];
    end
    always @(spike_out_source_array[507]) begin 
        spike_out_source507 = spike_out_source_array[507];
    end
    always @(spike_out_source_array[508]) begin 
        spike_out_source508 = spike_out_source_array[508];
    end
    always @(spike_out_source_array[509]) begin 
        spike_out_source509 = spike_out_source_array[509];
    end
    always @(spike_out_source_array[510]) begin 
        spike_out_source510 = spike_out_source_array[510];
    end
    always @(spike_out_source_array[511]) begin 
        spike_out_source511 = spike_out_source_array[511];
    end
    always @(spike_out_source_array[512]) begin 
        spike_out_source512 = spike_out_source_array[512];
    end
    always @(spike_out_source_array[513]) begin 
        spike_out_source513 = spike_out_source_array[513];
    end
    always @(spike_out_source_array[514]) begin 
        spike_out_source514 = spike_out_source_array[514];
    end
    always @(spike_out_source_array[515]) begin 
        spike_out_source515 = spike_out_source_array[515];
    end
    always @(spike_out_source_array[516]) begin 
        spike_out_source516 = spike_out_source_array[516];
    end
    always @(spike_out_source_array[517]) begin 
        spike_out_source517 = spike_out_source_array[517];
    end
    always @(spike_out_source_array[518]) begin 
        spike_out_source518 = spike_out_source_array[518];
    end
    always @(spike_out_source_array[519]) begin 
        spike_out_source519 = spike_out_source_array[519];
    end
    always @(spike_out_source_array[520]) begin 
        spike_out_source520 = spike_out_source_array[520];
    end
    always @(spike_out_source_array[521]) begin 
        spike_out_source521 = spike_out_source_array[521];
    end
    always @(spike_out_source_array[522]) begin 
        spike_out_source522 = spike_out_source_array[522];
    end
    always @(spike_out_source_array[523]) begin 
        spike_out_source523 = spike_out_source_array[523];
    end
    always @(spike_out_source_array[524]) begin 
        spike_out_source524 = spike_out_source_array[524];
    end
    always @(spike_out_source_array[525]) begin 
        spike_out_source525 = spike_out_source_array[525];
    end
    always @(spike_out_source_array[526]) begin 
        spike_out_source526 = spike_out_source_array[526];
    end
    always @(spike_out_source_array[527]) begin 
        spike_out_source527 = spike_out_source_array[527];
    end
    always @(spike_out_source_array[528]) begin 
        spike_out_source528 = spike_out_source_array[528];
    end
    always @(spike_out_source_array[529]) begin 
        spike_out_source529 = spike_out_source_array[529];
    end
    always @(spike_out_source_array[530]) begin 
        spike_out_source530 = spike_out_source_array[530];
    end
    always @(spike_out_source_array[531]) begin 
        spike_out_source531 = spike_out_source_array[531];
    end
    always @(spike_out_source_array[532]) begin 
        spike_out_source532 = spike_out_source_array[532];
    end
    always @(spike_out_source_array[533]) begin 
        spike_out_source533 = spike_out_source_array[533];
    end
    always @(spike_out_source_array[534]) begin 
        spike_out_source534 = spike_out_source_array[534];
    end
    always @(spike_out_source_array[535]) begin 
        spike_out_source535 = spike_out_source_array[535];
    end
    always @(spike_out_source_array[536]) begin 
        spike_out_source536 = spike_out_source_array[536];
    end
    always @(spike_out_source_array[537]) begin 
        spike_out_source537 = spike_out_source_array[537];
    end
    always @(spike_out_source_array[538]) begin 
        spike_out_source538 = spike_out_source_array[538];
    end
    always @(spike_out_source_array[539]) begin 
        spike_out_source539 = spike_out_source_array[539];
    end
    always @(spike_out_source_array[540]) begin 
        spike_out_source540 = spike_out_source_array[540];
    end
    always @(spike_out_source_array[541]) begin 
        spike_out_source541 = spike_out_source_array[541];
    end
    always @(spike_out_source_array[542]) begin 
        spike_out_source542 = spike_out_source_array[542];
    end
    always @(spike_out_source_array[543]) begin 
        spike_out_source543 = spike_out_source_array[543];
    end
    always @(spike_out_source_array[544]) begin 
        spike_out_source544 = spike_out_source_array[544];
    end
    always @(spike_out_source_array[545]) begin 
        spike_out_source545 = spike_out_source_array[545];
    end
    always @(spike_out_source_array[546]) begin 
        spike_out_source546 = spike_out_source_array[546];
    end
    always @(spike_out_source_array[547]) begin 
        spike_out_source547 = spike_out_source_array[547];
    end
    always @(spike_out_source_array[548]) begin 
        spike_out_source548 = spike_out_source_array[548];
    end
    always @(spike_out_source_array[549]) begin 
        spike_out_source549 = spike_out_source_array[549];
    end
    always @(spike_out_source_array[550]) begin 
        spike_out_source550 = spike_out_source_array[550];
    end
    always @(spike_out_source_array[551]) begin 
        spike_out_source551 = spike_out_source_array[551];
    end
    always @(spike_out_source_array[552]) begin 
        spike_out_source552 = spike_out_source_array[552];
    end
    always @(spike_out_source_array[553]) begin 
        spike_out_source553 = spike_out_source_array[553];
    end
    always @(spike_out_source_array[554]) begin 
        spike_out_source554 = spike_out_source_array[554];
    end
    always @(spike_out_source_array[555]) begin 
        spike_out_source555 = spike_out_source_array[555];
    end
    always @(spike_out_source_array[556]) begin 
        spike_out_source556 = spike_out_source_array[556];
    end
    always @(spike_out_source_array[557]) begin 
        spike_out_source557 = spike_out_source_array[557];
    end
    always @(spike_out_source_array[558]) begin 
        spike_out_source558 = spike_out_source_array[558];
    end
    always @(spike_out_source_array[559]) begin 
        spike_out_source559 = spike_out_source_array[559];
    end
    always @(spike_out_source_array[560]) begin 
        spike_out_source560 = spike_out_source_array[560];
    end
    always @(spike_out_source_array[561]) begin 
        spike_out_source561 = spike_out_source_array[561];
    end
    always @(spike_out_source_array[562]) begin 
        spike_out_source562 = spike_out_source_array[562];
    end
    always @(spike_out_source_array[563]) begin 
        spike_out_source563 = spike_out_source_array[563];
    end
    always @(spike_out_source_array[564]) begin 
        spike_out_source564 = spike_out_source_array[564];
    end
    always @(spike_out_source_array[565]) begin 
        spike_out_source565 = spike_out_source_array[565];
    end
    always @(spike_out_source_array[566]) begin 
        spike_out_source566 = spike_out_source_array[566];
    end
    always @(spike_out_source_array[567]) begin 
        spike_out_source567 = spike_out_source_array[567];
    end
    always @(spike_out_source_array[568]) begin 
        spike_out_source568 = spike_out_source_array[568];
    end
    always @(spike_out_source_array[569]) begin 
        spike_out_source569 = spike_out_source_array[569];
    end
    always @(spike_out_source_array[570]) begin 
        spike_out_source570 = spike_out_source_array[570];
    end
    always @(spike_out_source_array[571]) begin 
        spike_out_source571 = spike_out_source_array[571];
    end
    always @(spike_out_source_array[572]) begin 
        spike_out_source572 = spike_out_source_array[572];
    end
    always @(spike_out_source_array[573]) begin 
        spike_out_source573 = spike_out_source_array[573];
    end
    always @(spike_out_source_array[574]) begin 
        spike_out_source574 = spike_out_source_array[574];
    end
    always @(spike_out_source_array[575]) begin 
        spike_out_source575 = spike_out_source_array[575];
    end
    always @(spike_out_source_array[576]) begin 
        spike_out_source576 = spike_out_source_array[576];
    end
    always @(spike_out_source_array[577]) begin 
        spike_out_source577 = spike_out_source_array[577];
    end
    always @(spike_out_source_array[578]) begin 
        spike_out_source578 = spike_out_source_array[578];
    end
    always @(spike_out_source_array[579]) begin 
        spike_out_source579 = spike_out_source_array[579];
    end
    always @(spike_out_source_array[580]) begin 
        spike_out_source580 = spike_out_source_array[580];
    end
    always @(spike_out_source_array[581]) begin 
        spike_out_source581 = spike_out_source_array[581];
    end
    always @(spike_out_source_array[582]) begin 
        spike_out_source582 = spike_out_source_array[582];
    end
    always @(spike_out_source_array[583]) begin 
        spike_out_source583 = spike_out_source_array[583];
    end
    always @(spike_out_source_array[584]) begin 
        spike_out_source584 = spike_out_source_array[584];
    end
    always @(spike_out_source_array[585]) begin 
        spike_out_source585 = spike_out_source_array[585];
    end
    always @(spike_out_source_array[586]) begin 
        spike_out_source586 = spike_out_source_array[586];
    end
    always @(spike_out_source_array[587]) begin 
        spike_out_source587 = spike_out_source_array[587];
    end
    always @(spike_out_source_array[588]) begin 
        spike_out_source588 = spike_out_source_array[588];
    end
    always @(spike_out_source_array[589]) begin 
        spike_out_source589 = spike_out_source_array[589];
    end
    always @(spike_out_source_array[590]) begin 
        spike_out_source590 = spike_out_source_array[590];
    end
    always @(spike_out_source_array[591]) begin 
        spike_out_source591 = spike_out_source_array[591];
    end
    always @(spike_out_source_array[592]) begin 
        spike_out_source592 = spike_out_source_array[592];
    end
    always @(spike_out_source_array[593]) begin 
        spike_out_source593 = spike_out_source_array[593];
    end
    always @(spike_out_source_array[594]) begin 
        spike_out_source594 = spike_out_source_array[594];
    end
    always @(spike_out_source_array[595]) begin 
        spike_out_source595 = spike_out_source_array[595];
    end
    always @(spike_out_source_array[596]) begin 
        spike_out_source596 = spike_out_source_array[596];
    end
    always @(spike_out_source_array[597]) begin 
        spike_out_source597 = spike_out_source_array[597];
    end
    always @(spike_out_source_array[598]) begin 
        spike_out_source598 = spike_out_source_array[598];
    end
    always @(spike_out_source_array[599]) begin 
        spike_out_source599 = spike_out_source_array[599];
    end
    always @(spike_out_source_array[600]) begin 
        spike_out_source600 = spike_out_source_array[600];
    end
    always @(spike_out_source_array[601]) begin 
        spike_out_source601 = spike_out_source_array[601];
    end
    always @(spike_out_source_array[602]) begin 
        spike_out_source602 = spike_out_source_array[602];
    end
    always @(spike_out_source_array[603]) begin 
        spike_out_source603 = spike_out_source_array[603];
    end
    always @(spike_out_source_array[604]) begin 
        spike_out_source604 = spike_out_source_array[604];
    end
    always @(spike_out_source_array[605]) begin 
        spike_out_source605 = spike_out_source_array[605];
    end
    always @(spike_out_source_array[606]) begin 
        spike_out_source606 = spike_out_source_array[606];
    end
    always @(spike_out_source_array[607]) begin 
        spike_out_source607 = spike_out_source_array[607];
    end
    always @(spike_out_source_array[608]) begin 
        spike_out_source608 = spike_out_source_array[608];
    end
    always @(spike_out_source_array[609]) begin 
        spike_out_source609 = spike_out_source_array[609];
    end
    always @(spike_out_source_array[610]) begin 
        spike_out_source610 = spike_out_source_array[610];
    end
    always @(spike_out_source_array[611]) begin 
        spike_out_source611 = spike_out_source_array[611];
    end
    always @(spike_out_source_array[612]) begin 
        spike_out_source612 = spike_out_source_array[612];
    end
    always @(spike_out_source_array[613]) begin 
        spike_out_source613 = spike_out_source_array[613];
    end
    always @(spike_out_source_array[614]) begin 
        spike_out_source614 = spike_out_source_array[614];
    end
    always @(spike_out_source_array[615]) begin 
        spike_out_source615 = spike_out_source_array[615];
    end
    always @(spike_out_source_array[616]) begin 
        spike_out_source616 = spike_out_source_array[616];
    end
    always @(spike_out_source_array[617]) begin 
        spike_out_source617 = spike_out_source_array[617];
    end
    always @(spike_out_source_array[618]) begin 
        spike_out_source618 = spike_out_source_array[618];
    end
    always @(spike_out_source_array[619]) begin 
        spike_out_source619 = spike_out_source_array[619];
    end
    always @(spike_out_source_array[620]) begin 
        spike_out_source620 = spike_out_source_array[620];
    end
    always @(spike_out_source_array[621]) begin 
        spike_out_source621 = spike_out_source_array[621];
    end
    always @(spike_out_source_array[622]) begin 
        spike_out_source622 = spike_out_source_array[622];
    end
    always @(spike_out_source_array[623]) begin 
        spike_out_source623 = spike_out_source_array[623];
    end
    always @(spike_out_source_array[624]) begin 
        spike_out_source624 = spike_out_source_array[624];
    end
    always @(spike_out_source_array[625]) begin 
        spike_out_source625 = spike_out_source_array[625];
    end
    always @(spike_out_source_array[626]) begin 
        spike_out_source626 = spike_out_source_array[626];
    end
    always @(spike_out_source_array[627]) begin 
        spike_out_source627 = spike_out_source_array[627];
    end
    always @(spike_out_source_array[628]) begin 
        spike_out_source628 = spike_out_source_array[628];
    end
    always @(spike_out_source_array[629]) begin 
        spike_out_source629 = spike_out_source_array[629];
    end
    always @(spike_out_source_array[630]) begin 
        spike_out_source630 = spike_out_source_array[630];
    end
    always @(spike_out_source_array[631]) begin 
        spike_out_source631 = spike_out_source_array[631];
    end
    always @(spike_out_source_array[632]) begin 
        spike_out_source632 = spike_out_source_array[632];
    end
    always @(spike_out_source_array[633]) begin 
        spike_out_source633 = spike_out_source_array[633];
    end
    always @(spike_out_source_array[634]) begin 
        spike_out_source634 = spike_out_source_array[634];
    end
    always @(spike_out_source_array[635]) begin 
        spike_out_source635 = spike_out_source_array[635];
    end
    always @(spike_out_source_array[636]) begin 
        spike_out_source636 = spike_out_source_array[636];
    end
    always @(spike_out_source_array[637]) begin 
        spike_out_source637 = spike_out_source_array[637];
    end
    always @(spike_out_source_array[638]) begin 
        spike_out_source638 = spike_out_source_array[638];
    end
    always @(spike_out_source_array[639]) begin 
        spike_out_source639 = spike_out_source_array[639];
    end
    always @(spike_out_source_array[640]) begin 
        spike_out_source640 = spike_out_source_array[640];
    end
    always @(spike_out_source_array[641]) begin 
        spike_out_source641 = spike_out_source_array[641];
    end
    always @(spike_out_source_array[642]) begin 
        spike_out_source642 = spike_out_source_array[642];
    end
    always @(spike_out_source_array[643]) begin 
        spike_out_source643 = spike_out_source_array[643];
    end
    always @(spike_out_source_array[644]) begin 
        spike_out_source644 = spike_out_source_array[644];
    end
    always @(spike_out_source_array[645]) begin 
        spike_out_source645 = spike_out_source_array[645];
    end
    always @(spike_out_source_array[646]) begin 
        spike_out_source646 = spike_out_source_array[646];
    end
    always @(spike_out_source_array[647]) begin 
        spike_out_source647 = spike_out_source_array[647];
    end
    always @(spike_out_source_array[648]) begin 
        spike_out_source648 = spike_out_source_array[648];
    end
    always @(spike_out_source_array[649]) begin 
        spike_out_source649 = spike_out_source_array[649];
    end
    always @(spike_out_source_array[650]) begin 
        spike_out_source650 = spike_out_source_array[650];
    end
    always @(spike_out_source_array[651]) begin 
        spike_out_source651 = spike_out_source_array[651];
    end
    always @(spike_out_source_array[652]) begin 
        spike_out_source652 = spike_out_source_array[652];
    end
    always @(spike_out_source_array[653]) begin 
        spike_out_source653 = spike_out_source_array[653];
    end
    always @(spike_out_source_array[654]) begin 
        spike_out_source654 = spike_out_source_array[654];
    end
    always @(spike_out_source_array[655]) begin 
        spike_out_source655 = spike_out_source_array[655];
    end
    always @(spike_out_source_array[656]) begin 
        spike_out_source656 = spike_out_source_array[656];
    end
    always @(spike_out_source_array[657]) begin 
        spike_out_source657 = spike_out_source_array[657];
    end
    always @(spike_out_source_array[658]) begin 
        spike_out_source658 = spike_out_source_array[658];
    end
    always @(spike_out_source_array[659]) begin 
        spike_out_source659 = spike_out_source_array[659];
    end
    always @(spike_out_source_array[660]) begin 
        spike_out_source660 = spike_out_source_array[660];
    end
    always @(spike_out_source_array[661]) begin 
        spike_out_source661 = spike_out_source_array[661];
    end
    always @(spike_out_source_array[662]) begin 
        spike_out_source662 = spike_out_source_array[662];
    end
    always @(spike_out_source_array[663]) begin 
        spike_out_source663 = spike_out_source_array[663];
    end
    always @(spike_out_source_array[664]) begin 
        spike_out_source664 = spike_out_source_array[664];
    end
    always @(spike_out_source_array[665]) begin 
        spike_out_source665 = spike_out_source_array[665];
    end
    always @(spike_out_source_array[666]) begin 
        spike_out_source666 = spike_out_source_array[666];
    end
    always @(spike_out_source_array[667]) begin 
        spike_out_source667 = spike_out_source_array[667];
    end
    always @(spike_out_source_array[668]) begin 
        spike_out_source668 = spike_out_source_array[668];
    end
    always @(spike_out_source_array[669]) begin 
        spike_out_source669 = spike_out_source_array[669];
    end
    always @(spike_out_source_array[670]) begin 
        spike_out_source670 = spike_out_source_array[670];
    end
    always @(spike_out_source_array[671]) begin 
        spike_out_source671 = spike_out_source_array[671];
    end
    always @(spike_out_source_array[672]) begin 
        spike_out_source672 = spike_out_source_array[672];
    end
    always @(spike_out_source_array[673]) begin 
        spike_out_source673 = spike_out_source_array[673];
    end
    always @(spike_out_source_array[674]) begin 
        spike_out_source674 = spike_out_source_array[674];
    end
    always @(spike_out_source_array[675]) begin 
        spike_out_source675 = spike_out_source_array[675];
    end
    always @(spike_out_source_array[676]) begin 
        spike_out_source676 = spike_out_source_array[676];
    end
    always @(spike_out_source_array[677]) begin 
        spike_out_source677 = spike_out_source_array[677];
    end
    always @(spike_out_source_array[678]) begin 
        spike_out_source678 = spike_out_source_array[678];
    end
    always @(spike_out_source_array[679]) begin 
        spike_out_source679 = spike_out_source_array[679];
    end
    always @(spike_out_source_array[680]) begin 
        spike_out_source680 = spike_out_source_array[680];
    end
    always @(spike_out_source_array[681]) begin 
        spike_out_source681 = spike_out_source_array[681];
    end
    always @(spike_out_source_array[682]) begin 
        spike_out_source682 = spike_out_source_array[682];
    end
    always @(spike_out_source_array[683]) begin 
        spike_out_source683 = spike_out_source_array[683];
    end
    always @(spike_out_source_array[684]) begin 
        spike_out_source684 = spike_out_source_array[684];
    end
    always @(spike_out_source_array[685]) begin 
        spike_out_source685 = spike_out_source_array[685];
    end
    always @(spike_out_source_array[686]) begin 
        spike_out_source686 = spike_out_source_array[686];
    end
    always @(spike_out_source_array[687]) begin 
        spike_out_source687 = spike_out_source_array[687];
    end
    always @(spike_out_source_array[688]) begin 
        spike_out_source688 = spike_out_source_array[688];
    end
    always @(spike_out_source_array[689]) begin 
        spike_out_source689 = spike_out_source_array[689];
    end
    always @(spike_out_source_array[690]) begin 
        spike_out_source690 = spike_out_source_array[690];
    end
    always @(spike_out_source_array[691]) begin 
        spike_out_source691 = spike_out_source_array[691];
    end
    always @(spike_out_source_array[692]) begin 
        spike_out_source692 = spike_out_source_array[692];
    end
    always @(spike_out_source_array[693]) begin 
        spike_out_source693 = spike_out_source_array[693];
    end
    always @(spike_out_source_array[694]) begin 
        spike_out_source694 = spike_out_source_array[694];
    end
    always @(spike_out_source_array[695]) begin 
        spike_out_source695 = spike_out_source_array[695];
    end
    always @(spike_out_source_array[696]) begin 
        spike_out_source696 = spike_out_source_array[696];
    end
    always @(spike_out_source_array[697]) begin 
        spike_out_source697 = spike_out_source_array[697];
    end
    always @(spike_out_source_array[698]) begin 
        spike_out_source698 = spike_out_source_array[698];
    end
    always @(spike_out_source_array[699]) begin 
        spike_out_source699 = spike_out_source_array[699];
    end
    always @(spike_out_source_array[700]) begin 
        spike_out_source700 = spike_out_source_array[700];
    end
    always @(spike_out_source_array[701]) begin 
        spike_out_source701 = spike_out_source_array[701];
    end
    always @(spike_out_source_array[702]) begin 
        spike_out_source702 = spike_out_source_array[702];
    end
    always @(spike_out_source_array[703]) begin 
        spike_out_source703 = spike_out_source_array[703];
    end
    always @(spike_out_source_array[704]) begin 
        spike_out_source704 = spike_out_source_array[704];
    end
    always @(spike_out_source_array[705]) begin 
        spike_out_source705 = spike_out_source_array[705];
    end
    always @(spike_out_source_array[706]) begin 
        spike_out_source706 = spike_out_source_array[706];
    end
    always @(spike_out_source_array[707]) begin 
        spike_out_source707 = spike_out_source_array[707];
    end
    always @(spike_out_source_array[708]) begin 
        spike_out_source708 = spike_out_source_array[708];
    end
    always @(spike_out_source_array[709]) begin 
        spike_out_source709 = spike_out_source_array[709];
    end
    always @(spike_out_source_array[710]) begin 
        spike_out_source710 = spike_out_source_array[710];
    end
    always @(spike_out_source_array[711]) begin 
        spike_out_source711 = spike_out_source_array[711];
    end
    always @(spike_out_source_array[712]) begin 
        spike_out_source712 = spike_out_source_array[712];
    end
    always @(spike_out_source_array[713]) begin 
        spike_out_source713 = spike_out_source_array[713];
    end
    always @(spike_out_source_array[714]) begin 
        spike_out_source714 = spike_out_source_array[714];
    end
    always @(spike_out_source_array[715]) begin 
        spike_out_source715 = spike_out_source_array[715];
    end
    always @(spike_out_source_array[716]) begin 
        spike_out_source716 = spike_out_source_array[716];
    end
    always @(spike_out_source_array[717]) begin 
        spike_out_source717 = spike_out_source_array[717];
    end
    always @(spike_out_source_array[718]) begin 
        spike_out_source718 = spike_out_source_array[718];
    end
    always @(spike_out_source_array[719]) begin 
        spike_out_source719 = spike_out_source_array[719];
    end
    always @(spike_out_source_array[720]) begin 
        spike_out_source720 = spike_out_source_array[720];
    end
    always @(spike_out_source_array[721]) begin 
        spike_out_source721 = spike_out_source_array[721];
    end
    always @(spike_out_source_array[722]) begin 
        spike_out_source722 = spike_out_source_array[722];
    end
    always @(spike_out_source_array[723]) begin 
        spike_out_source723 = spike_out_source_array[723];
    end
    always @(spike_out_source_array[724]) begin 
        spike_out_source724 = spike_out_source_array[724];
    end
    always @(spike_out_source_array[725]) begin 
        spike_out_source725 = spike_out_source_array[725];
    end
    always @(spike_out_source_array[726]) begin 
        spike_out_source726 = spike_out_source_array[726];
    end
    always @(spike_out_source_array[727]) begin 
        spike_out_source727 = spike_out_source_array[727];
    end
    always @(spike_out_source_array[728]) begin 
        spike_out_source728 = spike_out_source_array[728];
    end
    always @(spike_out_source_array[729]) begin 
        spike_out_source729 = spike_out_source_array[729];
    end
    always @(spike_out_source_array[730]) begin 
        spike_out_source730 = spike_out_source_array[730];
    end
    always @(spike_out_source_array[731]) begin 
        spike_out_source731 = spike_out_source_array[731];
    end
    always @(spike_out_source_array[732]) begin 
        spike_out_source732 = spike_out_source_array[732];
    end
    always @(spike_out_source_array[733]) begin 
        spike_out_source733 = spike_out_source_array[733];
    end
    always @(spike_out_source_array[734]) begin 
        spike_out_source734 = spike_out_source_array[734];
    end
    always @(spike_out_source_array[735]) begin 
        spike_out_source735 = spike_out_source_array[735];
    end
    always @(spike_out_source_array[736]) begin 
        spike_out_source736 = spike_out_source_array[736];
    end
    always @(spike_out_source_array[737]) begin 
        spike_out_source737 = spike_out_source_array[737];
    end
    always @(spike_out_source_array[738]) begin 
        spike_out_source738 = spike_out_source_array[738];
    end
    always @(spike_out_source_array[739]) begin 
        spike_out_source739 = spike_out_source_array[739];
    end
    always @(spike_out_source_array[740]) begin 
        spike_out_source740 = spike_out_source_array[740];
    end
    always @(spike_out_source_array[741]) begin 
        spike_out_source741 = spike_out_source_array[741];
    end
    always @(spike_out_source_array[742]) begin 
        spike_out_source742 = spike_out_source_array[742];
    end
    always @(spike_out_source_array[743]) begin 
        spike_out_source743 = spike_out_source_array[743];
    end
    always @(spike_out_source_array[744]) begin 
        spike_out_source744 = spike_out_source_array[744];
    end
    always @(spike_out_source_array[745]) begin 
        spike_out_source745 = spike_out_source_array[745];
    end
    always @(spike_out_source_array[746]) begin 
        spike_out_source746 = spike_out_source_array[746];
    end
    always @(spike_out_source_array[747]) begin 
        spike_out_source747 = spike_out_source_array[747];
    end
    always @(spike_out_source_array[748]) begin 
        spike_out_source748 = spike_out_source_array[748];
    end
    always @(spike_out_source_array[749]) begin 
        spike_out_source749 = spike_out_source_array[749];
    end
    always @(spike_out_source_array[750]) begin 
        spike_out_source750 = spike_out_source_array[750];
    end
    always @(spike_out_source_array[751]) begin 
        spike_out_source751 = spike_out_source_array[751];
    end
    always @(spike_out_source_array[752]) begin 
        spike_out_source752 = spike_out_source_array[752];
    end
    always @(spike_out_source_array[753]) begin 
        spike_out_source753 = spike_out_source_array[753];
    end
    always @(spike_out_source_array[754]) begin 
        spike_out_source754 = spike_out_source_array[754];
    end
    always @(spike_out_source_array[755]) begin 
        spike_out_source755 = spike_out_source_array[755];
    end
    always @(spike_out_source_array[756]) begin 
        spike_out_source756 = spike_out_source_array[756];
    end
    always @(spike_out_source_array[757]) begin 
        spike_out_source757 = spike_out_source_array[757];
    end
    always @(spike_out_source_array[758]) begin 
        spike_out_source758 = spike_out_source_array[758];
    end
    always @(spike_out_source_array[759]) begin 
        spike_out_source759 = spike_out_source_array[759];
    end
    always @(spike_out_source_array[760]) begin 
        spike_out_source760 = spike_out_source_array[760];
    end
    always @(spike_out_source_array[761]) begin 
        spike_out_source761 = spike_out_source_array[761];
    end
    always @(spike_out_source_array[762]) begin 
        spike_out_source762 = spike_out_source_array[762];
    end
    always @(spike_out_source_array[763]) begin 
        spike_out_source763 = spike_out_source_array[763];
    end
    always @(spike_out_source_array[764]) begin 
        spike_out_source764 = spike_out_source_array[764];
    end
    always @(spike_out_source_array[765]) begin 
        spike_out_source765 = spike_out_source_array[765];
    end
    always @(spike_out_source_array[766]) begin 
        spike_out_source766 = spike_out_source_array[766];
    end
    always @(spike_out_source_array[767]) begin 
        spike_out_source767 = spike_out_source_array[767];
    end
    always @(spike_out_source_array[768]) begin 
        spike_out_source768 = spike_out_source_array[768];
    end
    always @(spike_out_source_array[769]) begin 
        spike_out_source769 = spike_out_source_array[769];
    end
    always @(spike_out_source_array[770]) begin 
        spike_out_source770 = spike_out_source_array[770];
    end
    always @(spike_out_source_array[771]) begin 
        spike_out_source771 = spike_out_source_array[771];
    end
    always @(spike_out_source_array[772]) begin 
        spike_out_source772 = spike_out_source_array[772];
    end
    always @(spike_out_source_array[773]) begin 
        spike_out_source773 = spike_out_source_array[773];
    end
    always @(spike_out_source_array[774]) begin 
        spike_out_source774 = spike_out_source_array[774];
    end
    always @(spike_out_source_array[775]) begin 
        spike_out_source775 = spike_out_source_array[775];
    end
    always @(spike_out_source_array[776]) begin 
        spike_out_source776 = spike_out_source_array[776];
    end
    always @(spike_out_source_array[777]) begin 
        spike_out_source777 = spike_out_source_array[777];
    end
    always @(spike_out_source_array[778]) begin 
        spike_out_source778 = spike_out_source_array[778];
    end
    always @(spike_out_source_array[779]) begin 
        spike_out_source779 = spike_out_source_array[779];
    end
    always @(spike_out_source_array[780]) begin 
        spike_out_source780 = spike_out_source_array[780];
    end
    always @(spike_out_source_array[781]) begin 
        spike_out_source781 = spike_out_source_array[781];
    end
    always @(spike_out_source_array[782]) begin 
        spike_out_source782 = spike_out_source_array[782];
    end
    always @(spike_out_source_array[783]) begin 
        spike_out_source783 = spike_out_source_array[783];
    end
    always @(spike_out_source_array[784]) begin 
        spike_out_source784 = spike_out_source_array[784];
    end
    always @(spike_out_source_array[785]) begin 
        spike_out_source785 = spike_out_source_array[785];
    end
    always @(spike_out_source_array[786]) begin 
        spike_out_source786 = spike_out_source_array[786];
    end
    always @(spike_out_source_array[787]) begin 
        spike_out_source787 = spike_out_source_array[787];
    end
    always @(spike_out_source_array[788]) begin 
        spike_out_source788 = spike_out_source_array[788];
    end
    always @(spike_out_source_array[789]) begin 
        spike_out_source789 = spike_out_source_array[789];
    end
    always @(spike_out_source_array[790]) begin 
        spike_out_source790 = spike_out_source_array[790];
    end
    always @(spike_out_source_array[791]) begin 
        spike_out_source791 = spike_out_source_array[791];
    end
    always @(spike_out_source_array[792]) begin 
        spike_out_source792 = spike_out_source_array[792];
    end
    always @(spike_out_source_array[793]) begin 
        spike_out_source793 = spike_out_source_array[793];
    end
    always @(spike_out_source_array[794]) begin 
        spike_out_source794 = spike_out_source_array[794];
    end
    always @(spike_out_source_array[795]) begin 
        spike_out_source795 = spike_out_source_array[795];
    end
    always @(spike_out_source_array[796]) begin 
        spike_out_source796 = spike_out_source_array[796];
    end
    always @(spike_out_source_array[797]) begin 
        spike_out_source797 = spike_out_source_array[797];
    end
    always @(spike_out_source_array[798]) begin 
        spike_out_source798 = spike_out_source_array[798];
    end
    always @(spike_out_source_array[799]) begin 
        spike_out_source799 = spike_out_source_array[799];
    end
    always @(spike_out_source_array[800]) begin 
        spike_out_source800 = spike_out_source_array[800];
    end
    always @(spike_out_source_array[801]) begin 
        spike_out_source801 = spike_out_source_array[801];
    end
    always @(spike_out_source_array[802]) begin 
        spike_out_source802 = spike_out_source_array[802];
    end
    always @(spike_out_source_array[803]) begin 
        spike_out_source803 = spike_out_source_array[803];
    end
    always @(spike_out_source_array[804]) begin 
        spike_out_source804 = spike_out_source_array[804];
    end
    always @(spike_out_source_array[805]) begin 
        spike_out_source805 = spike_out_source_array[805];
    end
    always @(spike_out_source_array[806]) begin 
        spike_out_source806 = spike_out_source_array[806];
    end
    always @(spike_out_source_array[807]) begin 
        spike_out_source807 = spike_out_source_array[807];
    end
    always @(spike_out_source_array[808]) begin 
        spike_out_source808 = spike_out_source_array[808];
    end
    always @(spike_out_source_array[809]) begin 
        spike_out_source809 = spike_out_source_array[809];
    end
    always @(spike_out_source_array[810]) begin 
        spike_out_source810 = spike_out_source_array[810];
    end
    always @(spike_out_source_array[811]) begin 
        spike_out_source811 = spike_out_source_array[811];
    end
    always @(spike_out_source_array[812]) begin 
        spike_out_source812 = spike_out_source_array[812];
    end
    always @(spike_out_source_array[813]) begin 
        spike_out_source813 = spike_out_source_array[813];
    end
    always @(spike_out_source_array[814]) begin 
        spike_out_source814 = spike_out_source_array[814];
    end
    always @(spike_out_source_array[815]) begin 
        spike_out_source815 = spike_out_source_array[815];
    end
    always @(spike_out_source_array[816]) begin 
        spike_out_source816 = spike_out_source_array[816];
    end
    always @(spike_out_source_array[817]) begin 
        spike_out_source817 = spike_out_source_array[817];
    end
    always @(spike_out_source_array[818]) begin 
        spike_out_source818 = spike_out_source_array[818];
    end
    always @(spike_out_source_array[819]) begin 
        spike_out_source819 = spike_out_source_array[819];
    end
    always @(spike_out_source_array[820]) begin 
        spike_out_source820 = spike_out_source_array[820];
    end
    always @(spike_out_source_array[821]) begin 
        spike_out_source821 = spike_out_source_array[821];
    end
    always @(spike_out_source_array[822]) begin 
        spike_out_source822 = spike_out_source_array[822];
    end
    always @(spike_out_source_array[823]) begin 
        spike_out_source823 = spike_out_source_array[823];
    end
    always @(spike_out_source_array[824]) begin 
        spike_out_source824 = spike_out_source_array[824];
    end
    always @(spike_out_source_array[825]) begin 
        spike_out_source825 = spike_out_source_array[825];
    end
    always @(spike_out_source_array[826]) begin 
        spike_out_source826 = spike_out_source_array[826];
    end
    always @(spike_out_source_array[827]) begin 
        spike_out_source827 = spike_out_source_array[827];
    end
    always @(spike_out_source_array[828]) begin 
        spike_out_source828 = spike_out_source_array[828];
    end
    always @(spike_out_source_array[829]) begin 
        spike_out_source829 = spike_out_source_array[829];
    end
    always @(spike_out_source_array[830]) begin 
        spike_out_source830 = spike_out_source_array[830];
    end
    always @(spike_out_source_array[831]) begin 
        spike_out_source831 = spike_out_source_array[831];
    end
    always @(spike_out_source_array[832]) begin 
        spike_out_source832 = spike_out_source_array[832];
    end
    always @(spike_out_source_array[833]) begin 
        spike_out_source833 = spike_out_source_array[833];
    end
    always @(spike_out_source_array[834]) begin 
        spike_out_source834 = spike_out_source_array[834];
    end
    always @(spike_out_source_array[835]) begin 
        spike_out_source835 = spike_out_source_array[835];
    end
    always @(spike_out_source_array[836]) begin 
        spike_out_source836 = spike_out_source_array[836];
    end
    always @(spike_out_source_array[837]) begin 
        spike_out_source837 = spike_out_source_array[837];
    end
    always @(spike_out_source_array[838]) begin 
        spike_out_source838 = spike_out_source_array[838];
    end
    always @(spike_out_source_array[839]) begin 
        spike_out_source839 = spike_out_source_array[839];
    end
    always @(spike_out_source_array[840]) begin 
        spike_out_source840 = spike_out_source_array[840];
    end
    always @(spike_out_source_array[841]) begin 
        spike_out_source841 = spike_out_source_array[841];
    end
    always @(spike_out_source_array[842]) begin 
        spike_out_source842 = spike_out_source_array[842];
    end
    always @(spike_out_source_array[843]) begin 
        spike_out_source843 = spike_out_source_array[843];
    end
    always @(spike_out_source_array[844]) begin 
        spike_out_source844 = spike_out_source_array[844];
    end
    always @(spike_out_source_array[845]) begin 
        spike_out_source845 = spike_out_source_array[845];
    end
    always @(spike_out_source_array[846]) begin 
        spike_out_source846 = spike_out_source_array[846];
    end
    always @(spike_out_source_array[847]) begin 
        spike_out_source847 = spike_out_source_array[847];
    end
    always @(spike_out_source_array[848]) begin 
        spike_out_source848 = spike_out_source_array[848];
    end
    always @(spike_out_source_array[849]) begin 
        spike_out_source849 = spike_out_source_array[849];
    end
    always @(spike_out_source_array[850]) begin 
        spike_out_source850 = spike_out_source_array[850];
    end
    always @(spike_out_source_array[851]) begin 
        spike_out_source851 = spike_out_source_array[851];
    end
    always @(spike_out_source_array[852]) begin 
        spike_out_source852 = spike_out_source_array[852];
    end
    always @(spike_out_source_array[853]) begin 
        spike_out_source853 = spike_out_source_array[853];
    end
    always @(spike_out_source_array[854]) begin 
        spike_out_source854 = spike_out_source_array[854];
    end
    always @(spike_out_source_array[855]) begin 
        spike_out_source855 = spike_out_source_array[855];
    end
    always @(spike_out_source_array[856]) begin 
        spike_out_source856 = spike_out_source_array[856];
    end
    always @(spike_out_source_array[857]) begin 
        spike_out_source857 = spike_out_source_array[857];
    end
    always @(spike_out_source_array[858]) begin 
        spike_out_source858 = spike_out_source_array[858];
    end
    always @(spike_out_source_array[859]) begin 
        spike_out_source859 = spike_out_source_array[859];
    end
    always @(spike_out_source_array[860]) begin 
        spike_out_source860 = spike_out_source_array[860];
    end
    always @(spike_out_source_array[861]) begin 
        spike_out_source861 = spike_out_source_array[861];
    end
    always @(spike_out_source_array[862]) begin 
        spike_out_source862 = spike_out_source_array[862];
    end
    always @(spike_out_source_array[863]) begin 
        spike_out_source863 = spike_out_source_array[863];
    end
    always @(spike_out_source_array[864]) begin 
        spike_out_source864 = spike_out_source_array[864];
    end
    always @(spike_out_source_array[865]) begin 
        spike_out_source865 = spike_out_source_array[865];
    end
    always @(spike_out_source_array[866]) begin 
        spike_out_source866 = spike_out_source_array[866];
    end
    always @(spike_out_source_array[867]) begin 
        spike_out_source867 = spike_out_source_array[867];
    end
    always @(spike_out_source_array[868]) begin 
        spike_out_source868 = spike_out_source_array[868];
    end
    always @(spike_out_source_array[869]) begin 
        spike_out_source869 = spike_out_source_array[869];
    end
    always @(spike_out_source_array[870]) begin 
        spike_out_source870 = spike_out_source_array[870];
    end
    always @(spike_out_source_array[871]) begin 
        spike_out_source871 = spike_out_source_array[871];
    end
    always @(spike_out_source_array[872]) begin 
        spike_out_source872 = spike_out_source_array[872];
    end
    always @(spike_out_source_array[873]) begin 
        spike_out_source873 = spike_out_source_array[873];
    end
    always @(spike_out_source_array[874]) begin 
        spike_out_source874 = spike_out_source_array[874];
    end
    always @(spike_out_source_array[875]) begin 
        spike_out_source875 = spike_out_source_array[875];
    end
    always @(spike_out_source_array[876]) begin 
        spike_out_source876 = spike_out_source_array[876];
    end
    always @(spike_out_source_array[877]) begin 
        spike_out_source877 = spike_out_source_array[877];
    end
    always @(spike_out_source_array[878]) begin 
        spike_out_source878 = spike_out_source_array[878];
    end
    always @(spike_out_source_array[879]) begin 
        spike_out_source879 = spike_out_source_array[879];
    end
    always @(spike_out_source_array[880]) begin 
        spike_out_source880 = spike_out_source_array[880];
    end
    always @(spike_out_source_array[881]) begin 
        spike_out_source881 = spike_out_source_array[881];
    end
    always @(spike_out_source_array[882]) begin 
        spike_out_source882 = spike_out_source_array[882];
    end
    always @(spike_out_source_array[883]) begin 
        spike_out_source883 = spike_out_source_array[883];
    end
    always @(spike_out_source_array[884]) begin 
        spike_out_source884 = spike_out_source_array[884];
    end
    always @(spike_out_source_array[885]) begin 
        spike_out_source885 = spike_out_source_array[885];
    end
    always @(spike_out_source_array[886]) begin 
        spike_out_source886 = spike_out_source_array[886];
    end
    always @(spike_out_source_array[887]) begin 
        spike_out_source887 = spike_out_source_array[887];
    end
    always @(spike_out_source_array[888]) begin 
        spike_out_source888 = spike_out_source_array[888];
    end
    always @(spike_out_source_array[889]) begin 
        spike_out_source889 = spike_out_source_array[889];
    end
    always @(spike_out_source_array[890]) begin 
        spike_out_source890 = spike_out_source_array[890];
    end
    always @(spike_out_source_array[891]) begin 
        spike_out_source891 = spike_out_source_array[891];
    end
    always @(spike_out_source_array[892]) begin 
        spike_out_source892 = spike_out_source_array[892];
    end
    always @(spike_out_source_array[893]) begin 
        spike_out_source893 = spike_out_source_array[893];
    end
    always @(spike_out_source_array[894]) begin 
        spike_out_source894 = spike_out_source_array[894];
    end
    always @(spike_out_source_array[895]) begin 
        spike_out_source895 = spike_out_source_array[895];
    end
    always @(spike_out_source_array[896]) begin 
        spike_out_source896 = spike_out_source_array[896];
    end
    always @(spike_out_source_array[897]) begin 
        spike_out_source897 = spike_out_source_array[897];
    end
    always @(spike_out_source_array[898]) begin 
        spike_out_source898 = spike_out_source_array[898];
    end
    always @(spike_out_source_array[899]) begin 
        spike_out_source899 = spike_out_source_array[899];
    end
    always @(spike_out_source_array[900]) begin 
        spike_out_source900 = spike_out_source_array[900];
    end
    always @(spike_out_source_array[901]) begin 
        spike_out_source901 = spike_out_source_array[901];
    end
    always @(spike_out_source_array[902]) begin 
        spike_out_source902 = spike_out_source_array[902];
    end
    always @(spike_out_source_array[903]) begin 
        spike_out_source903 = spike_out_source_array[903];
    end
    always @(spike_out_source_array[904]) begin 
        spike_out_source904 = spike_out_source_array[904];
    end
    always @(spike_out_source_array[905]) begin 
        spike_out_source905 = spike_out_source_array[905];
    end
    always @(spike_out_source_array[906]) begin 
        spike_out_source906 = spike_out_source_array[906];
    end
    always @(spike_out_source_array[907]) begin 
        spike_out_source907 = spike_out_source_array[907];
    end
    always @(spike_out_source_array[908]) begin 
        spike_out_source908 = spike_out_source_array[908];
    end
    always @(spike_out_source_array[909]) begin 
        spike_out_source909 = spike_out_source_array[909];
    end
    always @(spike_out_source_array[910]) begin 
        spike_out_source910 = spike_out_source_array[910];
    end
    always @(spike_out_source_array[911]) begin 
        spike_out_source911 = spike_out_source_array[911];
    end
    always @(spike_out_source_array[912]) begin 
        spike_out_source912 = spike_out_source_array[912];
    end
    always @(spike_out_source_array[913]) begin 
        spike_out_source913 = spike_out_source_array[913];
    end
    always @(spike_out_source_array[914]) begin 
        spike_out_source914 = spike_out_source_array[914];
    end
    always @(spike_out_source_array[915]) begin 
        spike_out_source915 = spike_out_source_array[915];
    end
    always @(spike_out_source_array[916]) begin 
        spike_out_source916 = spike_out_source_array[916];
    end
    always @(spike_out_source_array[917]) begin 
        spike_out_source917 = spike_out_source_array[917];
    end
    always @(spike_out_source_array[918]) begin 
        spike_out_source918 = spike_out_source_array[918];
    end
    always @(spike_out_source_array[919]) begin 
        spike_out_source919 = spike_out_source_array[919];
    end
    always @(spike_out_source_array[920]) begin 
        spike_out_source920 = spike_out_source_array[920];
    end
    always @(spike_out_source_array[921]) begin 
        spike_out_source921 = spike_out_source_array[921];
    end
    always @(spike_out_source_array[922]) begin 
        spike_out_source922 = spike_out_source_array[922];
    end
    always @(spike_out_source_array[923]) begin 
        spike_out_source923 = spike_out_source_array[923];
    end
    always @(spike_out_source_array[924]) begin 
        spike_out_source924 = spike_out_source_array[924];
    end
    always @(spike_out_source_array[925]) begin 
        spike_out_source925 = spike_out_source_array[925];
    end
    always @(spike_out_source_array[926]) begin 
        spike_out_source926 = spike_out_source_array[926];
    end
    always @(spike_out_source_array[927]) begin 
        spike_out_source927 = spike_out_source_array[927];
    end
    always @(spike_out_source_array[928]) begin 
        spike_out_source928 = spike_out_source_array[928];
    end
    always @(spike_out_source_array[929]) begin 
        spike_out_source929 = spike_out_source_array[929];
    end
    always @(spike_out_source_array[930]) begin 
        spike_out_source930 = spike_out_source_array[930];
    end
    always @(spike_out_source_array[931]) begin 
        spike_out_source931 = spike_out_source_array[931];
    end
    always @(spike_out_source_array[932]) begin 
        spike_out_source932 = spike_out_source_array[932];
    end
    always @(spike_out_source_array[933]) begin 
        spike_out_source933 = spike_out_source_array[933];
    end
    always @(spike_out_source_array[934]) begin 
        spike_out_source934 = spike_out_source_array[934];
    end
    always @(spike_out_source_array[935]) begin 
        spike_out_source935 = spike_out_source_array[935];
    end
    always @(spike_out_source_array[936]) begin 
        spike_out_source936 = spike_out_source_array[936];
    end
    always @(spike_out_source_array[937]) begin 
        spike_out_source937 = spike_out_source_array[937];
    end
    always @(spike_out_source_array[938]) begin 
        spike_out_source938 = spike_out_source_array[938];
    end
    always @(spike_out_source_array[939]) begin 
        spike_out_source939 = spike_out_source_array[939];
    end
    always @(spike_out_source_array[940]) begin 
        spike_out_source940 = spike_out_source_array[940];
    end
    always @(spike_out_source_array[941]) begin 
        spike_out_source941 = spike_out_source_array[941];
    end
    always @(spike_out_source_array[942]) begin 
        spike_out_source942 = spike_out_source_array[942];
    end
    always @(spike_out_source_array[943]) begin 
        spike_out_source943 = spike_out_source_array[943];
    end
    always @(spike_out_source_array[944]) begin 
        spike_out_source944 = spike_out_source_array[944];
    end
    always @(spike_out_source_array[945]) begin 
        spike_out_source945 = spike_out_source_array[945];
    end
    always @(spike_out_source_array[946]) begin 
        spike_out_source946 = spike_out_source_array[946];
    end
    always @(spike_out_source_array[947]) begin 
        spike_out_source947 = spike_out_source_array[947];
    end
    always @(spike_out_source_array[948]) begin 
        spike_out_source948 = spike_out_source_array[948];
    end
    always @(spike_out_source_array[949]) begin 
        spike_out_source949 = spike_out_source_array[949];
    end
    always @(spike_out_source_array[950]) begin 
        spike_out_source950 = spike_out_source_array[950];
    end
    always @(spike_out_source_array[951]) begin 
        spike_out_source951 = spike_out_source_array[951];
    end
    always @(spike_out_source_array[952]) begin 
        spike_out_source952 = spike_out_source_array[952];
    end
    always @(spike_out_source_array[953]) begin 
        spike_out_source953 = spike_out_source_array[953];
    end
    always @(spike_out_source_array[954]) begin 
        spike_out_source954 = spike_out_source_array[954];
    end
    always @(spike_out_source_array[955]) begin 
        spike_out_source955 = spike_out_source_array[955];
    end
    always @(spike_out_source_array[956]) begin 
        spike_out_source956 = spike_out_source_array[956];
    end
    always @(spike_out_source_array[957]) begin 
        spike_out_source957 = spike_out_source_array[957];
    end
    always @(spike_out_source_array[958]) begin 
        spike_out_source958 = spike_out_source_array[958];
    end
    always @(spike_out_source_array[959]) begin 
        spike_out_source959 = spike_out_source_array[959];
    end
    always @(spike_out_source_array[960]) begin 
        spike_out_source960 = spike_out_source_array[960];
    end
    always @(spike_out_source_array[961]) begin 
        spike_out_source961 = spike_out_source_array[961];
    end
    always @(spike_out_source_array[962]) begin 
        spike_out_source962 = spike_out_source_array[962];
    end
    always @(spike_out_source_array[963]) begin 
        spike_out_source963 = spike_out_source_array[963];
    end
    always @(spike_out_source_array[964]) begin 
        spike_out_source964 = spike_out_source_array[964];
    end
    always @(spike_out_source_array[965]) begin 
        spike_out_source965 = spike_out_source_array[965];
    end
    always @(spike_out_source_array[966]) begin 
        spike_out_source966 = spike_out_source_array[966];
    end
    always @(spike_out_source_array[967]) begin 
        spike_out_source967 = spike_out_source_array[967];
    end
    always @(spike_out_source_array[968]) begin 
        spike_out_source968 = spike_out_source_array[968];
    end
    always @(spike_out_source_array[969]) begin 
        spike_out_source969 = spike_out_source_array[969];
    end
    always @(spike_out_source_array[970]) begin 
        spike_out_source970 = spike_out_source_array[970];
    end
    always @(spike_out_source_array[971]) begin 
        spike_out_source971 = spike_out_source_array[971];
    end
    always @(spike_out_source_array[972]) begin 
        spike_out_source972 = spike_out_source_array[972];
    end
    always @(spike_out_source_array[973]) begin 
        spike_out_source973 = spike_out_source_array[973];
    end
    always @(spike_out_source_array[974]) begin 
        spike_out_source974 = spike_out_source_array[974];
    end
    always @(spike_out_source_array[975]) begin 
        spike_out_source975 = spike_out_source_array[975];
    end
    always @(spike_out_source_array[976]) begin 
        spike_out_source976 = spike_out_source_array[976];
    end
    always @(spike_out_source_array[977]) begin 
        spike_out_source977 = spike_out_source_array[977];
    end
    always @(spike_out_source_array[978]) begin 
        spike_out_source978 = spike_out_source_array[978];
    end
    always @(spike_out_source_array[979]) begin 
        spike_out_source979 = spike_out_source_array[979];
    end
    always @(spike_out_source_array[980]) begin 
        spike_out_source980 = spike_out_source_array[980];
    end
    always @(spike_out_source_array[981]) begin 
        spike_out_source981 = spike_out_source_array[981];
    end
    always @(spike_out_source_array[982]) begin 
        spike_out_source982 = spike_out_source_array[982];
    end
    always @(spike_out_source_array[983]) begin 
        spike_out_source983 = spike_out_source_array[983];
    end
    always @(spike_out_source_array[984]) begin 
        spike_out_source984 = spike_out_source_array[984];
    end
    always @(spike_out_source_array[985]) begin 
        spike_out_source985 = spike_out_source_array[985];
    end
    always @(spike_out_source_array[986]) begin 
        spike_out_source986 = spike_out_source_array[986];
    end
    always @(spike_out_source_array[987]) begin 
        spike_out_source987 = spike_out_source_array[987];
    end
    always @(spike_out_source_array[988]) begin 
        spike_out_source988 = spike_out_source_array[988];
    end
    always @(spike_out_source_array[989]) begin 
        spike_out_source989 = spike_out_source_array[989];
    end
    always @(spike_out_source_array[990]) begin 
        spike_out_source990 = spike_out_source_array[990];
    end
    always @(spike_out_source_array[991]) begin 
        spike_out_source991 = spike_out_source_array[991];
    end
    always @(spike_out_source_array[992]) begin 
        spike_out_source992 = spike_out_source_array[992];
    end
    always @(spike_out_source_array[993]) begin 
        spike_out_source993 = spike_out_source_array[993];
    end
    always @(spike_out_source_array[994]) begin 
        spike_out_source994 = spike_out_source_array[994];
    end
    always @(spike_out_source_array[995]) begin 
        spike_out_source995 = spike_out_source_array[995];
    end
    always @(spike_out_source_array[996]) begin 
        spike_out_source996 = spike_out_source_array[996];
    end
    always @(spike_out_source_array[997]) begin 
        spike_out_source997 = spike_out_source_array[997];
    end
    always @(spike_out_source_array[998]) begin 
        spike_out_source998 = spike_out_source_array[998];
    end
    always @(spike_out_source_array[999]) begin 
        spike_out_source999 = spike_out_source_array[999];
    end
    always @(spike_out_source_array[1000]) begin 
        spike_out_source1000 = spike_out_source_array[1000];
    end
    always @(spike_out_source_array[1001]) begin 
        spike_out_source1001 = spike_out_source_array[1001];
    end
    always @(spike_out_source_array[1002]) begin 
        spike_out_source1002 = spike_out_source_array[1002];
    end
    always @(spike_out_source_array[1003]) begin 
        spike_out_source1003 = spike_out_source_array[1003];
    end
    always @(spike_out_source_array[1004]) begin 
        spike_out_source1004 = spike_out_source_array[1004];
    end
    always @(spike_out_source_array[1005]) begin 
        spike_out_source1005 = spike_out_source_array[1005];
    end
    always @(spike_out_source_array[1006]) begin 
        spike_out_source1006 = spike_out_source_array[1006];
    end
    always @(spike_out_source_array[1007]) begin 
        spike_out_source1007 = spike_out_source_array[1007];
    end
    always @(spike_out_source_array[1008]) begin 
        spike_out_source1008 = spike_out_source_array[1008];
    end
    always @(spike_out_source_array[1009]) begin 
        spike_out_source1009 = spike_out_source_array[1009];
    end
    always @(spike_out_source_array[1010]) begin 
        spike_out_source1010 = spike_out_source_array[1010];
    end
    always @(spike_out_source_array[1011]) begin 
        spike_out_source1011 = spike_out_source_array[1011];
    end
    always @(spike_out_source_array[1012]) begin 
        spike_out_source1012 = spike_out_source_array[1012];
    end
    always @(spike_out_source_array[1013]) begin 
        spike_out_source1013 = spike_out_source_array[1013];
    end
    always @(spike_out_source_array[1014]) begin 
        spike_out_source1014 = spike_out_source_array[1014];
    end
    always @(spike_out_source_array[1015]) begin 
        spike_out_source1015 = spike_out_source_array[1015];
    end
    always @(spike_out_source_array[1016]) begin 
        spike_out_source1016 = spike_out_source_array[1016];
    end
    always @(spike_out_source_array[1017]) begin 
        spike_out_source1017 = spike_out_source_array[1017];
    end
    always @(spike_out_source_array[1018]) begin 
        spike_out_source1018 = spike_out_source_array[1018];
    end
    always @(spike_out_source_array[1019]) begin 
        spike_out_source1019 = spike_out_source_array[1019];
    end
    always @(spike_out_source_array[1020]) begin 
        spike_out_source1020 = spike_out_source_array[1020];
    end
    always @(spike_out_source_array[1021]) begin 
        spike_out_source1021 = spike_out_source_array[1021];
    end
    always @(spike_out_source_array[1022]) begin 
        spike_out_source1022 = spike_out_source_array[1022];
    end
    always @(spike_out_source_array[1023]) begin 
        spike_out_source1023 = spike_out_source_array[1023];
    end
    reg[18:0] i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21;
    reg[18:0] j1, j2, j3, j4, j5, j6, j7, j8, j9, j10, j11, j12, j13, j14, j15, j16, j17, j18, j19, j20, j21, module network_interface_scaled (
        input wire spike0,
    input wire spike1,    input wire spike2,    input wire spike3,    input wire spike4,    input wire spike5,    input wire spike6,    input wire spike7,    input wire spike8,    input wire spike9,    input wire spike10,    input wire spike11,    input wire spike12,    input wire spike13,    input wire spike14,    input wire spike15,    input wire spike16,    input wire spike17,    input wire spike18,    input wire spike19,    input wire spike20,    input wire spike21,    input wire spike22,    input wire spike23,    input wire spike24,    input wire spike25,    input wire spike26,    input wire spike27,    input wire spike28,    input wire spike29,    input wire spike30,    input wire spike31,    input wire spike32,    input wire spike33,    input wire spike34,    input wire spike35,    input wire spike36,    input wire spike37,    input wire spike38,    input wire spike39,    input wire spike40,    input wire spike41,    input wire spike42,    input wire spike43,    input wire spike44,    input wire spike45,    input wire spike46,    input wire spike47,    input wire spike48,    input wire spike49,    input wire spike50,    input wire spike51,    input wire spike52,    input wire spike53,    input wire spike54,    input wire spike55,    input wire spike56,    input wire spike57,    input wire spike58,    input wire spike59,    input wire spike60,    input wire spike61,    input wire spike62,    input wire spike63,    input wire spike64,    input wire spike65,    input wire spike66,    input wire spike67,    input wire spike68,    input wire spike69,    input wire spike70,    input wire spike71,    input wire spike72,    input wire spike73,    input wire spike74,    input wire spike75,    input wire spike76,    input wire spike77,    input wire spike78,    input wire spike79,    input wire spike80,    input wire spike81,    input wire spike82,    input wire spike83,    input wire spike84,    input wire spike85,    input wire spike86,    input wire spike87,    input wire spike88,    input wire spike89,    input wire spike90,    input wire spike91,    input wire spike92,    input wire spike93,    input wire spike94,    input wire spike95,    input wire spike96,    input wire spike97,    input wire spike98,    input wire spike99,    input wire spike100,
    input wire spike101,    input wire spike102,    input wire spike103,    input wire spike104,    input wire spike105,    input wire spike106,    input wire spike107,    input wire spike108,    input wire spike109,    input wire spike110,    input wire spike111,    input wire spike112,    input wire spike113,    input wire spike114,    input wire spike115,    input wire spike116,    input wire spike117,    input wire spike118,    input wire spike119,    input wire spike120,    input wire spike121,    input wire spike122,    input wire spike123,    input wire spike124,    input wire spike125,    input wire spike126,    input wire spike127,    input wire spike128,    input wire spike129,    input wire spike130,    input wire spike131,    input wire spike132,    input wire spike133,    input wire spike134,    input wire spike135,    input wire spike136,    input wire spike137,    input wire spike138,    input wire spike139,    input wire spike140,    input wire spike141,    input wire spike142,    input wire spike143,    input wire spike144,    input wire spike145,    input wire spike146,    input wire spike147,    input wire spike148,    input wire spike149,    input wire spike150,    input wire spike151,    input wire spike152,    input wire spike153,    input wire spike154,    input wire spike155,    input wire spike156,    input wire spike157,    input wire spike158,    input wire spike159,    input wire spike160,    input wire spike161,    input wire spike162,    input wire spike163,    input wire spike164,    input wire spike165,    input wire spike166,    input wire spike167,    input wire spike168,    input wire spike169,    input wire spike170,    input wire spike171,    input wire spike172,    input wire spike173,    input wire spike174,    input wire spike175,    input wire spike176,    input wire spike177,    input wire spike178,    input wire spike179,    input wire spike180,    input wire spike181,    input wire spike182,    input wire spike183,    input wire spike184,    input wire spike185,    input wire spike186,    input wire spike187,    input wire spike188,    input wire spike189,    input wire spike190,    input wire spike191,    input wire spike192,    input wire spike193,    input wire spike194,    input wire spike195,    input wire spike196,    input wire spike197,    input wire spike198,    input wire spike199,    input wire spike200,
    input wire spike201,    input wire spike202,    input wire spike203,    input wire spike204,    input wire spike205,    input wire spike206,    input wire spike207,    input wire spike208,    input wire spike209,    input wire spike210,    input wire spike211,    input wire spike212,    input wire spike213,    input wire spike214,    input wire spike215,    input wire spike216,    input wire spike217,    input wire spike218,    input wire spike219,    input wire spike220,    input wire spike221,    input wire spike222,    input wire spike223,    input wire spike224,    input wire spike225,    input wire spike226,    input wire spike227,    input wire spike228,    input wire spike229,    input wire spike230,    input wire spike231,    input wire spike232,    input wire spike233,    input wire spike234,    input wire spike235,    input wire spike236,    input wire spike237,    input wire spike238,    input wire spike239,    input wire spike240,    input wire spike241,    input wire spike242,    input wire spike243,    input wire spike244,    input wire spike245,    input wire spike246,    input wire spike247,    input wire spike248,    input wire spike249,    input wire spike250,    input wire spike251,    input wire spike252,    input wire spike253,    input wire spike254,    input wire spike255,    input wire spike256,    input wire spike257,    input wire spike258,    input wire spike259,    input wire spike260,    input wire spike261,    input wire spike262,    input wire spike263,    input wire spike264,    input wire spike265,    input wire spike266,    input wire spike267,    input wire spike268,    input wire spike269,    input wire spike270,    input wire spike271,    input wire spike272,    input wire spike273,    input wire spike274,    input wire spike275,    input wire spike276,    input wire spike277,    input wire spike278,    input wire spike279,    input wire spike280,    input wire spike281,    input wire spike282,    input wire spike283,    input wire spike284,    input wire spike285,    input wire spike286,    input wire spike287,    input wire spike288,    input wire spike289,    input wire spike290,    input wire spike291,    input wire spike292,    input wire spike293,    input wire spike294,    input wire spike295,    input wire spike296,    input wire spike297,    input wire spike298,    input wire spike299,    input wire spike300,
    input wire spike301,    input wire spike302,    input wire spike303,    input wire spike304,    input wire spike305,    input wire spike306,    input wire spike307,    input wire spike308,    input wire spike309,    input wire spike310,    input wire spike311,    input wire spike312,    input wire spike313,    input wire spike314,    input wire spike315,    input wire spike316,    input wire spike317,    input wire spike318,    input wire spike319,    input wire spike320,    input wire spike321,    input wire spike322,    input wire spike323,    input wire spike324,    input wire spike325,    input wire spike326,    input wire spike327,    input wire spike328,    input wire spike329,    input wire spike330,    input wire spike331,    input wire spike332,    input wire spike333,    input wire spike334,    input wire spike335,    input wire spike336,    input wire spike337,    input wire spike338,    input wire spike339,    input wire spike340,    input wire spike341,    input wire spike342,    input wire spike343,    input wire spike344,    input wire spike345,    input wire spike346,    input wire spike347,    input wire spike348,    input wire spike349,    input wire spike350,    input wire spike351,    input wire spike352,    input wire spike353,    input wire spike354,    input wire spike355,    input wire spike356,    input wire spike357,    input wire spike358,    input wire spike359,    input wire spike360,    input wire spike361,    input wire spike362,    input wire spike363,    input wire spike364,    input wire spike365,    input wire spike366,    input wire spike367,    input wire spike368,    input wire spike369,    input wire spike370,    input wire spike371,    input wire spike372,    input wire spike373,    input wire spike374,    input wire spike375,    input wire spike376,    input wire spike377,    input wire spike378,    input wire spike379,    input wire spike380,    input wire spike381,    input wire spike382,    input wire spike383,    input wire spike384,    input wire spike385,    input wire spike386,    input wire spike387,    input wire spike388,    input wire spike389,    input wire spike390,    input wire spike391,    input wire spike392,    input wire spike393,    input wire spike394,    input wire spike395,    input wire spike396,    input wire spike397,    input wire spike398,    input wire spike399,    input wire spike400,
    input wire spike401,    input wire spike402,    input wire spike403,    input wire spike404,    input wire spike405,    input wire spike406,    input wire spike407,    input wire spike408,    input wire spike409,    input wire spike410,    input wire spike411,    input wire spike412,    input wire spike413,    input wire spike414,    input wire spike415,    input wire spike416,    input wire spike417,    input wire spike418,    input wire spike419,    input wire spike420,    input wire spike421,    input wire spike422,    input wire spike423,    input wire spike424,    input wire spike425,    input wire spike426,    input wire spike427,    input wire spike428,    input wire spike429,    input wire spike430,    input wire spike431,    input wire spike432,    input wire spike433,    input wire spike434,    input wire spike435,    input wire spike436,    input wire spike437,    input wire spike438,    input wire spike439,    input wire spike440,    input wire spike441,    input wire spike442,    input wire spike443,    input wire spike444,    input wire spike445,    input wire spike446,    input wire spike447,    input wire spike448,    input wire spike449,    input wire spike450,    input wire spike451,    input wire spike452,    input wire spike453,    input wire spike454,    input wire spike455,    input wire spike456,    input wire spike457,    input wire spike458,    input wire spike459,    input wire spike460,    input wire spike461,    input wire spike462,    input wire spike463,    input wire spike464,    input wire spike465,    input wire spike466,    input wire spike467,    input wire spike468,    input wire spike469,    input wire spike470,    input wire spike471,    input wire spike472,    input wire spike473,    input wire spike474,    input wire spike475,    input wire spike476,    input wire spike477,    input wire spike478,    input wire spike479,    input wire spike480,    input wire spike481,    input wire spike482,    input wire spike483,    input wire spike484,    input wire spike485,    input wire spike486,    input wire spike487,    input wire spike488,    input wire spike489,    input wire spike490,    input wire spike491,    input wire spike492,    input wire spike493,    input wire spike494,    input wire spike495,    input wire spike496,    input wire spike497,    input wire spike498,    input wire spike499,    input wire spike500,
    input wire spike501,    input wire spike502,    input wire spike503,    input wire spike504,    input wire spike505,    input wire spike506,    input wire spike507,    input wire spike508,    input wire spike509,    input wire spike510,    input wire spike511,    input wire spike512,    input wire spike513,    input wire spike514,    input wire spike515,    input wire spike516,    input wire spike517,    input wire spike518,    input wire spike519,    input wire spike520,    input wire spike521,    input wire spike522,    input wire spike523,    input wire spike524,    input wire spike525,    input wire spike526,    input wire spike527,    input wire spike528,    input wire spike529,    input wire spike530,    input wire spike531,    input wire spike532,    input wire spike533,    input wire spike534,    input wire spike535,    input wire spike536,    input wire spike537,    input wire spike538,    input wire spike539,    input wire spike540,    input wire spike541,    input wire spike542,    input wire spike543,    input wire spike544,    input wire spike545,    input wire spike546,    input wire spike547,    input wire spike548,    input wire spike549,    input wire spike550,    input wire spike551,    input wire spike552,    input wire spike553,    input wire spike554,    input wire spike555,    input wire spike556,    input wire spike557,    input wire spike558,    input wire spike559,    input wire spike560,    input wire spike561,    input wire spike562,    input wire spike563,    input wire spike564,    input wire spike565,    input wire spike566,    input wire spike567,    input wire spike568,    input wire spike569,    input wire spike570,    input wire spike571,    input wire spike572,    input wire spike573,    input wire spike574,    input wire spike575,    input wire spike576,    input wire spike577,    input wire spike578,    input wire spike579,    input wire spike580,    input wire spike581,    input wire spike582,    input wire spike583,    input wire spike584,    input wire spike585,    input wire spike586,    input wire spike587,    input wire spike588,    input wire spike589,    input wire spike590,    input wire spike591,    input wire spike592,    input wire spike593,    input wire spike594,    input wire spike595,    input wire spike596,    input wire spike597,    input wire spike598,    input wire spike599,    input wire spike600,
    input wire spike601,    input wire spike602,    input wire spike603,    input wire spike604,    input wire spike605,    input wire spike606,    input wire spike607,    input wire spike608,    input wire spike609,    input wire spike610,    input wire spike611,    input wire spike612,    input wire spike613,    input wire spike614,    input wire spike615,    input wire spike616,    input wire spike617,    input wire spike618,    input wire spike619,    input wire spike620,    input wire spike621,    input wire spike622,    input wire spike623,    input wire spike624,    input wire spike625,    input wire spike626,    input wire spike627,    input wire spike628,    input wire spike629,    input wire spike630,    input wire spike631,    input wire spike632,    input wire spike633,    input wire spike634,    input wire spike635,    input wire spike636,    input wire spike637,    input wire spike638,    input wire spike639,    input wire spike640,    input wire spike641,    input wire spike642,    input wire spike643,    input wire spike644,    input wire spike645,    input wire spike646,    input wire spike647,    input wire spike648,    input wire spike649,    input wire spike650,    input wire spike651,    input wire spike652,    input wire spike653,    input wire spike654,    input wire spike655,    input wire spike656,    input wire spike657,    input wire spike658,    input wire spike659,    input wire spike660,    input wire spike661,    input wire spike662,    input wire spike663,    input wire spike664,    input wire spike665,    input wire spike666,    input wire spike667,    input wire spike668,    input wire spike669,    input wire spike670,    input wire spike671,    input wire spike672,    input wire spike673,    input wire spike674,    input wire spike675,    input wire spike676,    input wire spike677,    input wire spike678,    input wire spike679,    input wire spike680,    input wire spike681,    input wire spike682,    input wire spike683,    input wire spike684,    input wire spike685,    input wire spike686,    input wire spike687,    input wire spike688,    input wire spike689,    input wire spike690,    input wire spike691,    input wire spike692,    input wire spike693,    input wire spike694,    input wire spike695,    input wire spike696,    input wire spike697,    input wire spike698,    input wire spike699,    input wire spike700,
    input wire spike701,    input wire spike702,    input wire spike703,    input wire spike704,    input wire spike705,    input wire spike706,    input wire spike707,    input wire spike708,    input wire spike709,    input wire spike710,    input wire spike711,    input wire spike712,    input wire spike713,    input wire spike714,    input wire spike715,    input wire spike716,    input wire spike717,    input wire spike718,    input wire spike719,    input wire spike720,    input wire spike721,    input wire spike722,    input wire spike723,    input wire spike724,    input wire spike725,    input wire spike726,    input wire spike727,    input wire spike728,    input wire spike729,    input wire spike730,    input wire spike731,    input wire spike732,    input wire spike733,    input wire spike734,    input wire spike735,    input wire spike736,    input wire spike737,    input wire spike738,    input wire spike739,    input wire spike740,    input wire spike741,    input wire spike742,    input wire spike743,    input wire spike744,    input wire spike745,    input wire spike746,    input wire spike747,    input wire spike748,    input wire spike749,    input wire spike750,    input wire spike751,    input wire spike752,    input wire spike753,    input wire spike754,    input wire spike755,    input wire spike756,    input wire spike757,    input wire spike758,    input wire spike759,    input wire spike760,    input wire spike761,    input wire spike762,    input wire spike763,    input wire spike764,    input wire spike765,    input wire spike766,    input wire spike767,    input wire spike768,    input wire spike769,    input wire spike770,    input wire spike771,    input wire spike772,    input wire spike773,    input wire spike774,    input wire spike775,    input wire spike776,    input wire spike777,    input wire spike778,    input wire spike779,    input wire spike780,    input wire spike781,    input wire spike782,    input wire spike783,    input wire spike784,    input wire spike785,    input wire spike786,    input wire spike787,    input wire spike788,    input wire spike789,    input wire spike790,    input wire spike791,    input wire spike792,    input wire spike793,    input wire spike794,    input wire spike795,    input wire spike796,    input wire spike797,    input wire spike798,    input wire spike799,    input wire spike800,
    input wire spike801,    input wire spike802,    input wire spike803,    input wire spike804,    input wire spike805,    input wire spike806,    input wire spike807,    input wire spike808,    input wire spike809,    input wire spike810,    input wire spike811,    input wire spike812,    input wire spike813,    input wire spike814,    input wire spike815,    input wire spike816,    input wire spike817,    input wire spike818,    input wire spike819,    input wire spike820,    input wire spike821,    input wire spike822,    input wire spike823,    input wire spike824,    input wire spike825,    input wire spike826,    input wire spike827,    input wire spike828,    input wire spike829,    input wire spike830,    input wire spike831,    input wire spike832,    input wire spike833,    input wire spike834,    input wire spike835,    input wire spike836,    input wire spike837,    input wire spike838,    input wire spike839,    input wire spike840,    input wire spike841,    input wire spike842,    input wire spike843,    input wire spike844,    input wire spike845,    input wire spike846,    input wire spike847,    input wire spike848,    input wire spike849,    input wire spike850,    input wire spike851,    input wire spike852,    input wire spike853,    input wire spike854,    input wire spike855,    input wire spike856,    input wire spike857,    input wire spike858,    input wire spike859,    input wire spike860,    input wire spike861,    input wire spike862,    input wire spike863,    input wire spike864,    input wire spike865,    input wire spike866,    input wire spike867,    input wire spike868,    input wire spike869,    input wire spike870,    input wire spike871,    input wire spike872,    input wire spike873,    input wire spike874,    input wire spike875,    input wire spike876,    input wire spike877,    input wire spike878,    input wire spike879,    input wire spike880,    input wire spike881,    input wire spike882,    input wire spike883,    input wire spike884,    input wire spike885,    input wire spike886,    input wire spike887,    input wire spike888,    input wire spike889,    input wire spike890,    input wire spike891,    input wire spike892,    input wire spike893,    input wire spike894,    input wire spike895,    input wire spike896,    input wire spike897,    input wire spike898,    input wire spike899,    input wire spike900,
    input wire spike901,    input wire spike902,    input wire spike903,    input wire spike904,    input wire spike905,    input wire spike906,    input wire spike907,    input wire spike908,    input wire spike909,    input wire spike910,    input wire spike911,    input wire spike912,    input wire spike913,    input wire spike914,    input wire spike915,    input wire spike916,    input wire spike917,    input wire spike918,    input wire spike919,    input wire spike920,    input wire spike921,    input wire spike922,    input wire spike923,    input wire spike924,    input wire spike925,    input wire spike926,    input wire spike927,    input wire spike928,    input wire spike929,    input wire spike930,    input wire spike931,    input wire spike932,    input wire spike933,    input wire spike934,    input wire spike935,    input wire spike936,    input wire spike937,    input wire spike938,    input wire spike939,    input wire spike940,    input wire spike941,    input wire spike942,    input wire spike943,    input wire spike944,    input wire spike945,    input wire spike946,    input wire spike947,    input wire spike948,    input wire spike949,    input wire spike950,    input wire spike951,    input wire spike952,    input wire spike953,    input wire spike954,    input wire spike955,    input wire spike956,    input wire spike957,    input wire spike958,    input wire spike959,    input wire spike960,    input wire spike961,    input wire spike962,    input wire spike963,    input wire spike964,    input wire spike965,    input wire spike966,    input wire spike967,    input wire spike968,    input wire spike969,    input wire spike970,    input wire spike971,    input wire spike972,    input wire spike973,    input wire spike974,    input wire spike975,    input wire spike976,    input wire spike977,    input wire spike978,    input wire spike979,    input wire spike980,    input wire spike981,    input wire spike982,    input wire spike983,    input wire spike984,    input wire spike985,    input wire spike986,    input wire spike987,    input wire spike988,    input wire spike989,    input wire spike990,    input wire spike991,    input wire spike992,    input wire spike993,    input wire spike994,    input wire spike995,    input wire spike996,    input wire spike997,    input wire spike998,    input wire spike999,    input wire spike1000,
    input wire spike1001,    input wire spike1002,    input wire spike1003,    input wire spike1004,    input wire spike1005,    input wire spike1006,    input wire spike1007,    input wire spike1008,    input wire spike1009,    input wire spike1010,    input wire spike1011,    input wire spike1012,    input wire spike1013,    input wire spike1014,    input wire spike1015,    input wire spike1016,    input wire spike1017,    input wire spike1018,    input wire spike1019,    input wire spike1020,    input wire spike1021,    input wire spike1022,    input wire spike1023,
output reg[11:0]     spike_out_source0,
    spike_out_source1,    spike_out_source2,    spike_out_source3,    spike_out_source4,    spike_out_source5,    spike_out_source6,    spike_out_source7,    spike_out_source8,    spike_out_source9,    spike_out_source10,    spike_out_source11,    spike_out_source12,    spike_out_source13,    spike_out_source14,    spike_out_source15,    spike_out_source16,    spike_out_source17,    spike_out_source18,    spike_out_source19,    spike_out_source20,    spike_out_source21,    spike_out_source22,    spike_out_source23,    spike_out_source24,    spike_out_source25,    spike_out_source26,    spike_out_source27,    spike_out_source28,    spike_out_source29,    spike_out_source30,    spike_out_source31,    spike_out_source32,    spike_out_source33,    spike_out_source34,    spike_out_source35,    spike_out_source36,    spike_out_source37,    spike_out_source38,    spike_out_source39,    spike_out_source40,    spike_out_source41,    spike_out_source42,    spike_out_source43,    spike_out_source44,    spike_out_source45,    spike_out_source46,    spike_out_source47,    spike_out_source48,    spike_out_source49,    spike_out_source50,    spike_out_source51,    spike_out_source52,    spike_out_source53,    spike_out_source54,    spike_out_source55,    spike_out_source56,    spike_out_source57,    spike_out_source58,    spike_out_source59,    spike_out_source60,    spike_out_source61,    spike_out_source62,    spike_out_source63,    spike_out_source64,    spike_out_source65,    spike_out_source66,    spike_out_source67,    spike_out_source68,    spike_out_source69,    spike_out_source70,    spike_out_source71,    spike_out_source72,    spike_out_source73,    spike_out_source74,    spike_out_source75,    spike_out_source76,    spike_out_source77,    spike_out_source78,    spike_out_source79,    spike_out_source80,    spike_out_source81,    spike_out_source82,    spike_out_source83,    spike_out_source84,    spike_out_source85,    spike_out_source86,    spike_out_source87,    spike_out_source88,    spike_out_source89,    spike_out_source90,    spike_out_source91,    spike_out_source92,    spike_out_source93,    spike_out_source94,    spike_out_source95,    spike_out_source96,    spike_out_source97,    spike_out_source98,    spike_out_source99,    spike_out_source100,
    spike_out_source101,    spike_out_source102,    spike_out_source103,    spike_out_source104,    spike_out_source105,    spike_out_source106,    spike_out_source107,    spike_out_source108,    spike_out_source109,    spike_out_source110,    spike_out_source111,    spike_out_source112,    spike_out_source113,    spike_out_source114,    spike_out_source115,    spike_out_source116,    spike_out_source117,    spike_out_source118,    spike_out_source119,    spike_out_source120,    spike_out_source121,    spike_out_source122,    spike_out_source123,    spike_out_source124,    spike_out_source125,    spike_out_source126,    spike_out_source127,    spike_out_source128,    spike_out_source129,    spike_out_source130,    spike_out_source131,    spike_out_source132,    spike_out_source133,    spike_out_source134,    spike_out_source135,    spike_out_source136,    spike_out_source137,    spike_out_source138,    spike_out_source139,    spike_out_source140,    spike_out_source141,    spike_out_source142,    spike_out_source143,    spike_out_source144,    spike_out_source145,    spike_out_source146,    spike_out_source147,    spike_out_source148,    spike_out_source149,    spike_out_source150,    spike_out_source151,    spike_out_source152,    spike_out_source153,    spike_out_source154,    spike_out_source155,    spike_out_source156,    spike_out_source157,    spike_out_source158,    spike_out_source159,    spike_out_source160,    spike_out_source161,    spike_out_source162,    spike_out_source163,    spike_out_source164,    spike_out_source165,    spike_out_source166,    spike_out_source167,    spike_out_source168,    spike_out_source169,    spike_out_source170,    spike_out_source171,    spike_out_source172,    spike_out_source173,    spike_out_source174,    spike_out_source175,    spike_out_source176,    spike_out_source177,    spike_out_source178,    spike_out_source179,    spike_out_source180,    spike_out_source181,    spike_out_source182,    spike_out_source183,    spike_out_source184,    spike_out_source185,    spike_out_source186,    spike_out_source187,    spike_out_source188,    spike_out_source189,    spike_out_source190,    spike_out_source191,    spike_out_source192,    spike_out_source193,    spike_out_source194,    spike_out_source195,    spike_out_source196,    spike_out_source197,    spike_out_source198,    spike_out_source199,    spike_out_source200,
    spike_out_source201,    spike_out_source202,    spike_out_source203,    spike_out_source204,    spike_out_source205,    spike_out_source206,    spike_out_source207,    spike_out_source208,    spike_out_source209,    spike_out_source210,    spike_out_source211,    spike_out_source212,    spike_out_source213,    spike_out_source214,    spike_out_source215,    spike_out_source216,    spike_out_source217,    spike_out_source218,    spike_out_source219,    spike_out_source220,    spike_out_source221,    spike_out_source222,    spike_out_source223,    spike_out_source224,    spike_out_source225,    spike_out_source226,    spike_out_source227,    spike_out_source228,    spike_out_source229,    spike_out_source230,    spike_out_source231,    spike_out_source232,    spike_out_source233,    spike_out_source234,    spike_out_source235,    spike_out_source236,    spike_out_source237,    spike_out_source238,    spike_out_source239,    spike_out_source240,    spike_out_source241,    spike_out_source242,    spike_out_source243,    spike_out_source244,    spike_out_source245,    spike_out_source246,    spike_out_source247,    spike_out_source248,    spike_out_source249,    spike_out_source250,    spike_out_source251,    spike_out_source252,    spike_out_source253,    spike_out_source254,    spike_out_source255,    spike_out_source256,    spike_out_source257,    spike_out_source258,    spike_out_source259,    spike_out_source260,    spike_out_source261,    spike_out_source262,    spike_out_source263,    spike_out_source264,    spike_out_source265,    spike_out_source266,    spike_out_source267,    spike_out_source268,    spike_out_source269,    spike_out_source270,    spike_out_source271,    spike_out_source272,    spike_out_source273,    spike_out_source274,    spike_out_source275,    spike_out_source276,    spike_out_source277,    spike_out_source278,    spike_out_source279,    spike_out_source280,    spike_out_source281,    spike_out_source282,    spike_out_source283,    spike_out_source284,    spike_out_source285,    spike_out_source286,    spike_out_source287,    spike_out_source288,    spike_out_source289,    spike_out_source290,    spike_out_source291,    spike_out_source292,    spike_out_source293,    spike_out_source294,    spike_out_source295,    spike_out_source296,    spike_out_source297,    spike_out_source298,    spike_out_source299,    spike_out_source300,
    spike_out_source301,    spike_out_source302,    spike_out_source303,    spike_out_source304,    spike_out_source305,    spike_out_source306,    spike_out_source307,    spike_out_source308,    spike_out_source309,    spike_out_source310,    spike_out_source311,    spike_out_source312,    spike_out_source313,    spike_out_source314,    spike_out_source315,    spike_out_source316,    spike_out_source317,    spike_out_source318,    spike_out_source319,    spike_out_source320,    spike_out_source321,    spike_out_source322,    spike_out_source323,    spike_out_source324,    spike_out_source325,    spike_out_source326,    spike_out_source327,    spike_out_source328,    spike_out_source329,    spike_out_source330,    spike_out_source331,    spike_out_source332,    spike_out_source333,    spike_out_source334,    spike_out_source335,    spike_out_source336,    spike_out_source337,    spike_out_source338,    spike_out_source339,    spike_out_source340,    spike_out_source341,    spike_out_source342,    spike_out_source343,    spike_out_source344,    spike_out_source345,    spike_out_source346,    spike_out_source347,    spike_out_source348,    spike_out_source349,    spike_out_source350,    spike_out_source351,    spike_out_source352,    spike_out_source353,    spike_out_source354,    spike_out_source355,    spike_out_source356,    spike_out_source357,    spike_out_source358,    spike_out_source359,    spike_out_source360,    spike_out_source361,    spike_out_source362,    spike_out_source363,    spike_out_source364,    spike_out_source365,    spike_out_source366,    spike_out_source367,    spike_out_source368,    spike_out_source369,    spike_out_source370,    spike_out_source371,    spike_out_source372,    spike_out_source373,    spike_out_source374,    spike_out_source375,    spike_out_source376,    spike_out_source377,    spike_out_source378,    spike_out_source379,    spike_out_source380,    spike_out_source381,    spike_out_source382,    spike_out_source383,    spike_out_source384,    spike_out_source385,    spike_out_source386,    spike_out_source387,    spike_out_source388,    spike_out_source389,    spike_out_source390,    spike_out_source391,    spike_out_source392,    spike_out_source393,    spike_out_source394,    spike_out_source395,    spike_out_source396,    spike_out_source397,    spike_out_source398,    spike_out_source399,    spike_out_source400,
    spike_out_source401,    spike_out_source402,    spike_out_source403,    spike_out_source404,    spike_out_source405,    spike_out_source406,    spike_out_source407,    spike_out_source408,    spike_out_source409,    spike_out_source410,    spike_out_source411,    spike_out_source412,    spike_out_source413,    spike_out_source414,    spike_out_source415,    spike_out_source416,    spike_out_source417,    spike_out_source418,    spike_out_source419,    spike_out_source420,    spike_out_source421,    spike_out_source422,    spike_out_source423,    spike_out_source424,    spike_out_source425,    spike_out_source426,    spike_out_source427,    spike_out_source428,    spike_out_source429,    spike_out_source430,    spike_out_source431,    spike_out_source432,    spike_out_source433,    spike_out_source434,    spike_out_source435,    spike_out_source436,    spike_out_source437,    spike_out_source438,    spike_out_source439,    spike_out_source440,    spike_out_source441,    spike_out_source442,    spike_out_source443,    spike_out_source444,    spike_out_source445,    spike_out_source446,    spike_out_source447,    spike_out_source448,    spike_out_source449,    spike_out_source450,    spike_out_source451,    spike_out_source452,    spike_out_source453,    spike_out_source454,    spike_out_source455,    spike_out_source456,    spike_out_source457,    spike_out_source458,    spike_out_source459,    spike_out_source460,    spike_out_source461,    spike_out_source462,    spike_out_source463,    spike_out_source464,    spike_out_source465,    spike_out_source466,    spike_out_source467,    spike_out_source468,    spike_out_source469,    spike_out_source470,    spike_out_source471,    spike_out_source472,    spike_out_source473,    spike_out_source474,    spike_out_source475,    spike_out_source476,    spike_out_source477,    spike_out_source478,    spike_out_source479,    spike_out_source480,    spike_out_source481,    spike_out_source482,    spike_out_source483,    spike_out_source484,    spike_out_source485,    spike_out_source486,    spike_out_source487,    spike_out_source488,    spike_out_source489,    spike_out_source490,    spike_out_source491,    spike_out_source492,    spike_out_source493,    spike_out_source494,    spike_out_source495,    spike_out_source496,    spike_out_source497,    spike_out_source498,    spike_out_source499,    spike_out_source500,
    spike_out_source501,    spike_out_source502,    spike_out_source503,    spike_out_source504,    spike_out_source505,    spike_out_source506,    spike_out_source507,    spike_out_source508,    spike_out_source509,    spike_out_source510,    spike_out_source511,    spike_out_source512,    spike_out_source513,    spike_out_source514,    spike_out_source515,    spike_out_source516,    spike_out_source517,    spike_out_source518,    spike_out_source519,    spike_out_source520,    spike_out_source521,    spike_out_source522,    spike_out_source523,    spike_out_source524,    spike_out_source525,    spike_out_source526,    spike_out_source527,    spike_out_source528,    spike_out_source529,    spike_out_source530,    spike_out_source531,    spike_out_source532,    spike_out_source533,    spike_out_source534,    spike_out_source535,    spike_out_source536,    spike_out_source537,    spike_out_source538,    spike_out_source539,    spike_out_source540,    spike_out_source541,    spike_out_source542,    spike_out_source543,    spike_out_source544,    spike_out_source545,    spike_out_source546,    spike_out_source547,    spike_out_source548,    spike_out_source549,    spike_out_source550,    spike_out_source551,    spike_out_source552,    spike_out_source553,    spike_out_source554,    spike_out_source555,    spike_out_source556,    spike_out_source557,    spike_out_source558,    spike_out_source559,    spike_out_source560,    spike_out_source561,    spike_out_source562,    spike_out_source563,    spike_out_source564,    spike_out_source565,    spike_out_source566,    spike_out_source567,    spike_out_source568,    spike_out_source569,    spike_out_source570,    spike_out_source571,    spike_out_source572,    spike_out_source573,    spike_out_source574,    spike_out_source575,    spike_out_source576,    spike_out_source577,    spike_out_source578,    spike_out_source579,    spike_out_source580,    spike_out_source581,    spike_out_source582,    spike_out_source583,    spike_out_source584,    spike_out_source585,    spike_out_source586,    spike_out_source587,    spike_out_source588,    spike_out_source589,    spike_out_source590,    spike_out_source591,    spike_out_source592,    spike_out_source593,    spike_out_source594,    spike_out_source595,    spike_out_source596,    spike_out_source597,    spike_out_source598,    spike_out_source599,    spike_out_source600,
    spike_out_source601,    spike_out_source602,    spike_out_source603,    spike_out_source604,    spike_out_source605,    spike_out_source606,    spike_out_source607,    spike_out_source608,    spike_out_source609,    spike_out_source610,    spike_out_source611,    spike_out_source612,    spike_out_source613,    spike_out_source614,    spike_out_source615,    spike_out_source616,    spike_out_source617,    spike_out_source618,    spike_out_source619,    spike_out_source620,    spike_out_source621,    spike_out_source622,    spike_out_source623,    spike_out_source624,    spike_out_source625,    spike_out_source626,    spike_out_source627,    spike_out_source628,    spike_out_source629,    spike_out_source630,    spike_out_source631,    spike_out_source632,    spike_out_source633,    spike_out_source634,    spike_out_source635,    spike_out_source636,    spike_out_source637,    spike_out_source638,    spike_out_source639,    spike_out_source640,    spike_out_source641,    spike_out_source642,    spike_out_source643,    spike_out_source644,    spike_out_source645,    spike_out_source646,    spike_out_source647,    spike_out_source648,    spike_out_source649,    spike_out_source650,    spike_out_source651,    spike_out_source652,    spike_out_source653,    spike_out_source654,    spike_out_source655,    spike_out_source656,    spike_out_source657,    spike_out_source658,    spike_out_source659,    spike_out_source660,    spike_out_source661,    spike_out_source662,    spike_out_source663,    spike_out_source664,    spike_out_source665,    spike_out_source666,    spike_out_source667,    spike_out_source668,    spike_out_source669,    spike_out_source670,    spike_out_source671,    spike_out_source672,    spike_out_source673,    spike_out_source674,    spike_out_source675,    spike_out_source676,    spike_out_source677,    spike_out_source678,    spike_out_source679,    spike_out_source680,    spike_out_source681,    spike_out_source682,    spike_out_source683,    spike_out_source684,    spike_out_source685,    spike_out_source686,    spike_out_source687,    spike_out_source688,    spike_out_source689,    spike_out_source690,    spike_out_source691,    spike_out_source692,    spike_out_source693,    spike_out_source694,    spike_out_source695,    spike_out_source696,    spike_out_source697,    spike_out_source698,    spike_out_source699,    spike_out_source700,
    spike_out_source701,    spike_out_source702,    spike_out_source703,    spike_out_source704,    spike_out_source705,    spike_out_source706,    spike_out_source707,    spike_out_source708,    spike_out_source709,    spike_out_source710,    spike_out_source711,    spike_out_source712,    spike_out_source713,    spike_out_source714,    spike_out_source715,    spike_out_source716,    spike_out_source717,    spike_out_source718,    spike_out_source719,    spike_out_source720,    spike_out_source721,    spike_out_source722,    spike_out_source723,    spike_out_source724,    spike_out_source725,    spike_out_source726,    spike_out_source727,    spike_out_source728,    spike_out_source729,    spike_out_source730,    spike_out_source731,    spike_out_source732,    spike_out_source733,    spike_out_source734,    spike_out_source735,    spike_out_source736,    spike_out_source737,    spike_out_source738,    spike_out_source739,    spike_out_source740,    spike_out_source741,    spike_out_source742,    spike_out_source743,    spike_out_source744,    spike_out_source745,    spike_out_source746,    spike_out_source747,    spike_out_source748,    spike_out_source749,    spike_out_source750,    spike_out_source751,    spike_out_source752,    spike_out_source753,    spike_out_source754,    spike_out_source755,    spike_out_source756,    spike_out_source757,    spike_out_source758,    spike_out_source759,    spike_out_source760,    spike_out_source761,    spike_out_source762,    spike_out_source763,    spike_out_source764,    spike_out_source765,    spike_out_source766,    spike_out_source767,    spike_out_source768,    spike_out_source769,    spike_out_source770,    spike_out_source771,    spike_out_source772,    spike_out_source773,    spike_out_source774,    spike_out_source775,    spike_out_source776,    spike_out_source777,    spike_out_source778,    spike_out_source779,    spike_out_source780,    spike_out_source781,    spike_out_source782,    spike_out_source783,    spike_out_source784,    spike_out_source785,    spike_out_source786,    spike_out_source787,    spike_out_source788,    spike_out_source789,    spike_out_source790,    spike_out_source791,    spike_out_source792,    spike_out_source793,    spike_out_source794,    spike_out_source795,    spike_out_source796,    spike_out_source797,    spike_out_source798,    spike_out_source799,    spike_out_source800,
    spike_out_source801,    spike_out_source802,    spike_out_source803,    spike_out_source804,    spike_out_source805,    spike_out_source806,    spike_out_source807,    spike_out_source808,    spike_out_source809,    spike_out_source810,    spike_out_source811,    spike_out_source812,    spike_out_source813,    spike_out_source814,    spike_out_source815,    spike_out_source816,    spike_out_source817,    spike_out_source818,    spike_out_source819,    spike_out_source820,    spike_out_source821,    spike_out_source822,    spike_out_source823,    spike_out_source824,    spike_out_source825,    spike_out_source826,    spike_out_source827,    spike_out_source828,    spike_out_source829,    spike_out_source830,    spike_out_source831,    spike_out_source832,    spike_out_source833,    spike_out_source834,    spike_out_source835,    spike_out_source836,    spike_out_source837,    spike_out_source838,    spike_out_source839,    spike_out_source840,    spike_out_source841,    spike_out_source842,    spike_out_source843,    spike_out_source844,    spike_out_source845,    spike_out_source846,    spike_out_source847,    spike_out_source848,    spike_out_source849,    spike_out_source850,    spike_out_source851,    spike_out_source852,    spike_out_source853,    spike_out_source854,    spike_out_source855,    spike_out_source856,    spike_out_source857,    spike_out_source858,    spike_out_source859,    spike_out_source860,    spike_out_source861,    spike_out_source862,    spike_out_source863,    spike_out_source864,    spike_out_source865,    spike_out_source866,    spike_out_source867,    spike_out_source868,    spike_out_source869,    spike_out_source870,    spike_out_source871,    spike_out_source872,    spike_out_source873,    spike_out_source874,    spike_out_source875,    spike_out_source876,    spike_out_source877,    spike_out_source878,    spike_out_source879,    spike_out_source880,    spike_out_source881,    spike_out_source882,    spike_out_source883,    spike_out_source884,    spike_out_source885,    spike_out_source886,    spike_out_source887,    spike_out_source888,    spike_out_source889,    spike_out_source890,    spike_out_source891,    spike_out_source892,    spike_out_source893,    spike_out_source894,    spike_out_source895,    spike_out_source896,    spike_out_source897,    spike_out_source898,    spike_out_source899,    spike_out_source900,
    spike_out_source901,    spike_out_source902,    spike_out_source903,    spike_out_source904,    spike_out_source905,    spike_out_source906,    spike_out_source907,    spike_out_source908,    spike_out_source909,    spike_out_source910,    spike_out_source911,    spike_out_source912,    spike_out_source913,    spike_out_source914,    spike_out_source915,    spike_out_source916,    spike_out_source917,    spike_out_source918,    spike_out_source919,    spike_out_source920,    spike_out_source921,    spike_out_source922,    spike_out_source923,    spike_out_source924,    spike_out_source925,    spike_out_source926,    spike_out_source927,    spike_out_source928,    spike_out_source929,    spike_out_source930,    spike_out_source931,    spike_out_source932,    spike_out_source933,    spike_out_source934,    spike_out_source935,    spike_out_source936,    spike_out_source937,    spike_out_source938,    spike_out_source939,    spike_out_source940,    spike_out_source941,    spike_out_source942,    spike_out_source943,    spike_out_source944,    spike_out_source945,    spike_out_source946,    spike_out_source947,    spike_out_source948,    spike_out_source949,    spike_out_source950,    spike_out_source951,    spike_out_source952,    spike_out_source953,    spike_out_source954,    spike_out_source955,    spike_out_source956,    spike_out_source957,    spike_out_source958,    spike_out_source959,    spike_out_source960,    spike_out_source961,    spike_out_source962,    spike_out_source963,    spike_out_source964,    spike_out_source965,    spike_out_source966,    spike_out_source967,    spike_out_source968,    spike_out_source969,    spike_out_source970,    spike_out_source971,    spike_out_source972,    spike_out_source973,    spike_out_source974,    spike_out_source975,    spike_out_source976,    spike_out_source977,    spike_out_source978,    spike_out_source979,    spike_out_source980,    spike_out_source981,    spike_out_source982,    spike_out_source983,    spike_out_source984,    spike_out_source985,    spike_out_source986,    spike_out_source987,    spike_out_source988,    spike_out_source989,    spike_out_source990,    spike_out_source991,    spike_out_source992,    spike_out_source993,    spike_out_source994,    spike_out_source995,    spike_out_source996,    spike_out_source997,    spike_out_source998,    spike_out_source999,    spike_out_source1000,
    spike_out_source1001,    spike_out_source1002,    spike_out_source1003,    spike_out_source1004,    spike_out_source1005,    spike_out_source1006,    spike_out_source1007,    spike_out_source1008,    spike_out_source1009,    spike_out_source1010,    spike_out_source1011,    spike_out_source1012,    spike_out_source1013,    spike_out_source1014,    spike_out_source1015,    spike_out_source1016,    spike_out_source1017,    spike_out_source1018,    spike_out_source1019,    spike_out_source1020,    spike_out_source1021,    spike_out_source1022,    spike_out_source1023,
    output wire output
);

    parameter number_of_neurons= 1024;
    reg spike_register[0:number_of_neurons-1];
    always @(clear, lock1, spike0, spike1, spike2, spike3, spike4, spike5, spike6, spike7, spike8, spike9, spike10, spike11, spike12, spike13, spike14, spike15, spike16, spike17, spike18, spike19, spike20, spike21, spike22, spike23, spike24, spike25, spike26, spike27, spike28, spike29, spike30, spike31, spike32, spike33, spike34, spike35, spike36, spike37, spike38, spike39, spike40, spike41, spike42, spike43, spike44, spike45, spike46, spike47, spike48, spike49) begin
        spike_register[0] = spike0;

        spike_register[1] = spike1;        spike_register[2] = spike2;        spike_register[3] = spike3;        spike_register[4] = spike4;        spike_register[5] = spike5;        spike_register[6] = spike6;        spike_register[7] = spike7;        spike_register[8] = spike8;        spike_register[9] = spike9;        spike_register[10] = spike10;        spike_register[11] = spike11;        spike_register[12] = spike12;        spike_register[13] = spike13;        spike_register[14] = spike14;        spike_register[15] = spike15;        spike_register[16] = spike16;        spike_register[17] = spike17;        spike_register[18] = spike18;        spike_register[19] = spike19;        spike_register[20] = spike20;        spike_register[21] = spike21;        spike_register[22] = spike22;        spike_register[23] = spike23;        spike_register[24] = spike24;        spike_register[25] = spike25;        spike_register[26] = spike26;        spike_register[27] = spike27;        spike_register[28] = spike28;        spike_register[29] = spike29;        spike_register[30] = spike30;        spike_register[31] = spike31;        spike_register[32] = spike32;        spike_register[33] = spike33;        spike_register[34] = spike34;        spike_register[35] = spike35;        spike_register[36] = spike36;        spike_register[37] = spike37;        spike_register[38] = spike38;        spike_register[39] = spike39;        spike_register[40] = spike40;        spike_register[41] = spike41;        spike_register[42] = spike42;        spike_register[43] = spike43;        spike_register[44] = spike44;        spike_register[45] = spike45;        spike_register[46] = spike46;        spike_register[47] = spike47;        spike_register[48] = spike48;        spike_register[49] = spike49;
        #0.5
        if(clear == 1'b0) begin
            for(i1 = 0; i1 <=49; i1= i1+1) begin
                if(spike_register[i1] == 1 && lock1 == 0) begin
                    lock1 = 1;
                    for(j1 = connection_pointer[i1]; j1 < connection_pointer[i1+1]; j1= j1+1) begin
                        packet1 = #0.1 {neuron_addresses[i1], downstream_connections[j1]};
                    end
                    spike_register[i1] = 0;
                    lock1 = 0;
                end
            end
        end

    end
    always @(clear, lock2, spike50, spike51, spike52, spike53, spike54, spike55, spike56, spike57, spike58, spike59, spike60, spike61, spike62, spike63, spike64, spike65, spike66, spike67, spike68, spike69, spike70, spike71, spike72, spike73, spike74, spike75, spike76, spike77, spike78, spike79, spike80, spike81, spike82, spike83, spike84, spike85, spike86, spike87, spike88, spike89, spike90, spike91, spike92, spike93, spike94, spike95, spike96, spike97, spike98, spike99) begin
        spike_register[50] = spike50;        spike_register[51] = spike51;        spike_register[52] = spike52;        spike_register[53] = spike53;        spike_register[54] = spike54;        spike_register[55] = spike55;        spike_register[56] = spike56;        spike_register[57] = spike57;        spike_register[58] = spike58;        spike_register[59] = spike59;        spike_register[60] = spike60;        spike_register[61] = spike61;        spike_register[62] = spike62;        spike_register[63] = spike63;        spike_register[64] = spike64;        spike_register[65] = spike65;        spike_register[66] = spike66;        spike_register[67] = spike67;        spike_register[68] = spike68;        spike_register[69] = spike69;        spike_register[70] = spike70;        spike_register[71] = spike71;        spike_register[72] = spike72;        spike_register[73] = spike73;        spike_register[74] = spike74;        spike_register[75] = spike75;        spike_register[76] = spike76;        spike_register[77] = spike77;        spike_register[78] = spike78;        spike_register[79] = spike79;        spike_register[80] = spike80;        spike_register[81] = spike81;        spike_register[82] = spike82;        spike_register[83] = spike83;        spike_register[84] = spike84;        spike_register[85] = spike85;        spike_register[86] = spike86;        spike_register[87] = spike87;        spike_register[88] = spike88;        spike_register[89] = spike89;        spike_register[90] = spike90;        spike_register[91] = spike91;        spike_register[92] = spike92;        spike_register[93] = spike93;        spike_register[94] = spike94;        spike_register[95] = spike95;        spike_register[96] = spike96;        spike_register[97] = spike97;        spike_register[98] = spike98;        spike_register[99] = spike99;
        #0.5
        if(clear == 1'b0) begin
            for(i2 = 50; i2 <=99; i2= i2+1) begin
                if(spike_register[i2] == 1 && lock2 == 0) begin
                    lock2 = 1;
                    for(j2 = connection_pointer[i2]; j2 < connection_pointer[i2+1]; j2= j2+1) begin
                        packet2 = #0.1 {neuron_addresses[i2], downstream_connections[j2]};
                    end
                    spike_register[i2] = 0;
                    lock2 = 0;
                end
            end
        end

    end
    always @(clear, lock3, spike100, spike101, spike102, spike103, spike104, spike105, spike106, spike107, spike108, spike109, spike110, spike111, spike112, spike113, spike114, spike115, spike116, spike117, spike118, spike119, spike120, spike121, spike122, spike123, spike124, spike125, spike126, spike127, spike128, spike129, spike130, spike131, spike132, spike133, spike134, spike135, spike136, spike137, spike138, spike139, spike140, spike141, spike142, spike143, spike144, spike145, spike146, spike147, spike148, spike149) begin
        spike_register[100] = spike100;

        spike_register[101] = spike101;        spike_register[102] = spike102;        spike_register[103] = spike103;        spike_register[104] = spike104;        spike_register[105] = spike105;        spike_register[106] = spike106;        spike_register[107] = spike107;        spike_register[108] = spike108;        spike_register[109] = spike109;        spike_register[110] = spike110;        spike_register[111] = spike111;        spike_register[112] = spike112;        spike_register[113] = spike113;        spike_register[114] = spike114;        spike_register[115] = spike115;        spike_register[116] = spike116;        spike_register[117] = spike117;        spike_register[118] = spike118;        spike_register[119] = spike119;        spike_register[120] = spike120;        spike_register[121] = spike121;        spike_register[122] = spike122;        spike_register[123] = spike123;        spike_register[124] = spike124;        spike_register[125] = spike125;        spike_register[126] = spike126;        spike_register[127] = spike127;        spike_register[128] = spike128;        spike_register[129] = spike129;        spike_register[130] = spike130;        spike_register[131] = spike131;        spike_register[132] = spike132;        spike_register[133] = spike133;        spike_register[134] = spike134;        spike_register[135] = spike135;        spike_register[136] = spike136;        spike_register[137] = spike137;        spike_register[138] = spike138;        spike_register[139] = spike139;        spike_register[140] = spike140;        spike_register[141] = spike141;        spike_register[142] = spike142;        spike_register[143] = spike143;        spike_register[144] = spike144;        spike_register[145] = spike145;        spike_register[146] = spike146;        spike_register[147] = spike147;        spike_register[148] = spike148;        spike_register[149] = spike149;
        #0.5
        if(clear == 1'b0) begin
            for(i3 = 100; i3 <=149; i3= i3+1) begin
                if(spike_register[i3] == 1 && lock3 == 0) begin
                    lock3 = 1;
                    for(j3 = connection_pointer[i3]; j3 < connection_pointer[i3+1]; j3= j3+1) begin
                        packet3 = #0.1 {neuron_addresses[i3], downstream_connections[j3]};
                    end
                    spike_register[i3] = 0;
                    lock3 = 0;
                end
            end
        end

    end
    always @(clear, lock4, spike150, spike151, spike152, spike153, spike154, spike155, spike156, spike157, spike158, spike159, spike160, spike161, spike162, spike163, spike164, spike165, spike166, spike167, spike168, spike169, spike170, spike171, spike172, spike173, spike174, spike175, spike176, spike177, spike178, spike179, spike180, spike181, spike182, spike183, spike184, spike185, spike186, spike187, spike188, spike189, spike190, spike191, spike192, spike193, spike194, spike195, spike196, spike197, spike198, spike199) begin
        spike_register[150] = spike150;        spike_register[151] = spike151;        spike_register[152] = spike152;        spike_register[153] = spike153;        spike_register[154] = spike154;        spike_register[155] = spike155;        spike_register[156] = spike156;        spike_register[157] = spike157;        spike_register[158] = spike158;        spike_register[159] = spike159;        spike_register[160] = spike160;        spike_register[161] = spike161;        spike_register[162] = spike162;        spike_register[163] = spike163;        spike_register[164] = spike164;        spike_register[165] = spike165;        spike_register[166] = spike166;        spike_register[167] = spike167;        spike_register[168] = spike168;        spike_register[169] = spike169;        spike_register[170] = spike170;        spike_register[171] = spike171;        spike_register[172] = spike172;        spike_register[173] = spike173;        spike_register[174] = spike174;        spike_register[175] = spike175;        spike_register[176] = spike176;        spike_register[177] = spike177;        spike_register[178] = spike178;        spike_register[179] = spike179;        spike_register[180] = spike180;        spike_register[181] = spike181;        spike_register[182] = spike182;        spike_register[183] = spike183;        spike_register[184] = spike184;        spike_register[185] = spike185;        spike_register[186] = spike186;        spike_register[187] = spike187;        spike_register[188] = spike188;        spike_register[189] = spike189;        spike_register[190] = spike190;        spike_register[191] = spike191;        spike_register[192] = spike192;        spike_register[193] = spike193;        spike_register[194] = spike194;        spike_register[195] = spike195;        spike_register[196] = spike196;        spike_register[197] = spike197;        spike_register[198] = spike198;        spike_register[199] = spike199;
        #0.5
        if(clear == 1'b0) begin
            for(i4 = 150; i4 <=199; i4= i4+1) begin
                if(spike_register[i4] == 1 && lock4 == 0) begin
                    lock4 = 1;
                    for(j4 = connection_pointer[i4]; j4 < connection_pointer[i4+1]; j4= j4+1) begin
                        packet4 = #0.1 {neuron_addresses[i4], downstream_connections[j4]};
                    end
                    spike_register[i4] = 0;
                    lock4 = 0;
                end
            end
        end

    end
    always @(clear, lock5, spike200, spike201, spike202, spike203, spike204, spike205, spike206, spike207, spike208, spike209, spike210, spike211, spike212, spike213, spike214, spike215, spike216, spike217, spike218, spike219, spike220, spike221, spike222, spike223, spike224, spike225, spike226, spike227, spike228, spike229, spike230, spike231, spike232, spike233, spike234, spike235, spike236, spike237, spike238, spike239, spike240, spike241, spike242, spike243, spike244, spike245, spike246, spike247, spike248, spike249) begin
        spike_register[200] = spike200;

        spike_register[201] = spike201;        spike_register[202] = spike202;        spike_register[203] = spike203;        spike_register[204] = spike204;        spike_register[205] = spike205;        spike_register[206] = spike206;        spike_register[207] = spike207;        spike_register[208] = spike208;        spike_register[209] = spike209;        spike_register[210] = spike210;        spike_register[211] = spike211;        spike_register[212] = spike212;        spike_register[213] = spike213;        spike_register[214] = spike214;        spike_register[215] = spike215;        spike_register[216] = spike216;        spike_register[217] = spike217;        spike_register[218] = spike218;        spike_register[219] = spike219;        spike_register[220] = spike220;        spike_register[221] = spike221;        spike_register[222] = spike222;        spike_register[223] = spike223;        spike_register[224] = spike224;        spike_register[225] = spike225;        spike_register[226] = spike226;        spike_register[227] = spike227;        spike_register[228] = spike228;        spike_register[229] = spike229;        spike_register[230] = spike230;        spike_register[231] = spike231;        spike_register[232] = spike232;        spike_register[233] = spike233;        spike_register[234] = spike234;        spike_register[235] = spike235;        spike_register[236] = spike236;        spike_register[237] = spike237;        spike_register[238] = spike238;        spike_register[239] = spike239;        spike_register[240] = spike240;        spike_register[241] = spike241;        spike_register[242] = spike242;        spike_register[243] = spike243;        spike_register[244] = spike244;        spike_register[245] = spike245;        spike_register[246] = spike246;        spike_register[247] = spike247;        spike_register[248] = spike248;        spike_register[249] = spike249;
        #0.5
        if(clear == 1'b0) begin
            for(i5 = 200; i5 <=249; i5= i5+1) begin
                if(spike_register[i5] == 1 && lock5 == 0) begin
                    lock5 = 1;
                    for(j5 = connection_pointer[i5]; j5 < connection_pointer[i5+1]; j5= j5+1) begin
                        packet5 = #0.1 {neuron_addresses[i5], downstream_connections[j5]};
                    end
                    spike_register[i5] = 0;
                    lock5 = 0;
                end
            end
        end

    end
    always @(clear, lock6, spike250, spike251, spike252, spike253, spike254, spike255, spike256, spike257, spike258, spike259, spike260, spike261, spike262, spike263, spike264, spike265, spike266, spike267, spike268, spike269, spike270, spike271, spike272, spike273, spike274, spike275, spike276, spike277, spike278, spike279, spike280, spike281, spike282, spike283, spike284, spike285, spike286, spike287, spike288, spike289, spike290, spike291, spike292, spike293, spike294, spike295, spike296, spike297, spike298, spike299) begin
        spike_register[250] = spike250;        spike_register[251] = spike251;        spike_register[252] = spike252;        spike_register[253] = spike253;        spike_register[254] = spike254;        spike_register[255] = spike255;        spike_register[256] = spike256;        spike_register[257] = spike257;        spike_register[258] = spike258;        spike_register[259] = spike259;        spike_register[260] = spike260;        spike_register[261] = spike261;        spike_register[262] = spike262;        spike_register[263] = spike263;        spike_register[264] = spike264;        spike_register[265] = spike265;        spike_register[266] = spike266;        spike_register[267] = spike267;        spike_register[268] = spike268;        spike_register[269] = spike269;        spike_register[270] = spike270;        spike_register[271] = spike271;        spike_register[272] = spike272;        spike_register[273] = spike273;        spike_register[274] = spike274;        spike_register[275] = spike275;        spike_register[276] = spike276;        spike_register[277] = spike277;        spike_register[278] = spike278;        spike_register[279] = spike279;        spike_register[280] = spike280;        spike_register[281] = spike281;        spike_register[282] = spike282;        spike_register[283] = spike283;        spike_register[284] = spike284;        spike_register[285] = spike285;        spike_register[286] = spike286;        spike_register[287] = spike287;        spike_register[288] = spike288;        spike_register[289] = spike289;        spike_register[290] = spike290;        spike_register[291] = spike291;        spike_register[292] = spike292;        spike_register[293] = spike293;        spike_register[294] = spike294;        spike_register[295] = spike295;        spike_register[296] = spike296;        spike_register[297] = spike297;        spike_register[298] = spike298;        spike_register[299] = spike299;
        #0.5
        if(clear == 1'b0) begin
            for(i6 = 250; i6 <=299; i6= i6+1) begin
                if(spike_register[i6] == 1 && lock6 == 0) begin
                    lock6 = 1;
                    for(j6 = connection_pointer[i6]; j6 < connection_pointer[i6+1]; j6= j6+1) begin
                        packet6 = #0.1 {neuron_addresses[i6], downstream_connections[j6]};
                    end
                    spike_register[i6] = 0;
                    lock6 = 0;
                end
            end
        end

    end
    always @(clear, lock7, spike300, spike301, spike302, spike303, spike304, spike305, spike306, spike307, spike308, spike309, spike310, spike311, spike312, spike313, spike314, spike315, spike316, spike317, spike318, spike319, spike320, spike321, spike322, spike323, spike324, spike325, spike326, spike327, spike328, spike329, spike330, spike331, spike332, spike333, spike334, spike335, spike336, spike337, spike338, spike339, spike340, spike341, spike342, spike343, spike344, spike345, spike346, spike347, spike348, spike349) begin
        spike_register[300] = spike300;

        spike_register[301] = spike301;        spike_register[302] = spike302;        spike_register[303] = spike303;        spike_register[304] = spike304;        spike_register[305] = spike305;        spike_register[306] = spike306;        spike_register[307] = spike307;        spike_register[308] = spike308;        spike_register[309] = spike309;        spike_register[310] = spike310;        spike_register[311] = spike311;        spike_register[312] = spike312;        spike_register[313] = spike313;        spike_register[314] = spike314;        spike_register[315] = spike315;        spike_register[316] = spike316;        spike_register[317] = spike317;        spike_register[318] = spike318;        spike_register[319] = spike319;        spike_register[320] = spike320;        spike_register[321] = spike321;        spike_register[322] = spike322;        spike_register[323] = spike323;        spike_register[324] = spike324;        spike_register[325] = spike325;        spike_register[326] = spike326;        spike_register[327] = spike327;        spike_register[328] = spike328;        spike_register[329] = spike329;        spike_register[330] = spike330;        spike_register[331] = spike331;        spike_register[332] = spike332;        spike_register[333] = spike333;        spike_register[334] = spike334;        spike_register[335] = spike335;        spike_register[336] = spike336;        spike_register[337] = spike337;        spike_register[338] = spike338;        spike_register[339] = spike339;        spike_register[340] = spike340;        spike_register[341] = spike341;        spike_register[342] = spike342;        spike_register[343] = spike343;        spike_register[344] = spike344;        spike_register[345] = spike345;        spike_register[346] = spike346;        spike_register[347] = spike347;        spike_register[348] = spike348;        spike_register[349] = spike349;
        #0.5
        if(clear == 1'b0) begin
            for(i7 = 300; i7 <=349; i7= i7+1) begin
                if(spike_register[i7] == 1 && lock7 == 0) begin
                    lock7 = 1;
                    for(j7 = connection_pointer[i7]; j7 < connection_pointer[i7+1]; j7= j7+1) begin
                        packet7 = #0.1 {neuron_addresses[i7], downstream_connections[j7]};
                    end
                    spike_register[i7] = 0;
                    lock7 = 0;
                end
            end
        end

    end
    always @(clear, lock8, spike350, spike351, spike352, spike353, spike354, spike355, spike356, spike357, spike358, spike359, spike360, spike361, spike362, spike363, spike364, spike365, spike366, spike367, spike368, spike369, spike370, spike371, spike372, spike373, spike374, spike375, spike376, spike377, spike378, spike379, spike380, spike381, spike382, spike383, spike384, spike385, spike386, spike387, spike388, spike389, spike390, spike391, spike392, spike393, spike394, spike395, spike396, spike397, spike398, spike399) begin
        spike_register[350] = spike350;        spike_register[351] = spike351;        spike_register[352] = spike352;        spike_register[353] = spike353;        spike_register[354] = spike354;        spike_register[355] = spike355;        spike_register[356] = spike356;        spike_register[357] = spike357;        spike_register[358] = spike358;        spike_register[359] = spike359;        spike_register[360] = spike360;        spike_register[361] = spike361;        spike_register[362] = spike362;        spike_register[363] = spike363;        spike_register[364] = spike364;        spike_register[365] = spike365;        spike_register[366] = spike366;        spike_register[367] = spike367;        spike_register[368] = spike368;        spike_register[369] = spike369;        spike_register[370] = spike370;        spike_register[371] = spike371;        spike_register[372] = spike372;        spike_register[373] = spike373;        spike_register[374] = spike374;        spike_register[375] = spike375;        spike_register[376] = spike376;        spike_register[377] = spike377;        spike_register[378] = spike378;        spike_register[379] = spike379;        spike_register[380] = spike380;        spike_register[381] = spike381;        spike_register[382] = spike382;        spike_register[383] = spike383;        spike_register[384] = spike384;        spike_register[385] = spike385;        spike_register[386] = spike386;        spike_register[387] = spike387;        spike_register[388] = spike388;        spike_register[389] = spike389;        spike_register[390] = spike390;        spike_register[391] = spike391;        spike_register[392] = spike392;        spike_register[393] = spike393;        spike_register[394] = spike394;        spike_register[395] = spike395;        spike_register[396] = spike396;        spike_register[397] = spike397;        spike_register[398] = spike398;        spike_register[399] = spike399;
        #0.5
        if(clear == 1'b0) begin
            for(i8 = 350; i8 <=399; i8= i8+1) begin
                if(spike_register[i8] == 1 && lock8 == 0) begin
                    lock8 = 1;
                    for(j8 = connection_pointer[i8]; j8 < connection_pointer[i8+1]; j8= j8+1) begin
                        packet8 = #0.1 {neuron_addresses[i8], downstream_connections[j8]};
                    end
                    spike_register[i8] = 0;
                    lock8 = 0;
                end
            end
        end

    end
    always @(clear, lock9, spike400, spike401, spike402, spike403, spike404, spike405, spike406, spike407, spike408, spike409, spike410, spike411, spike412, spike413, spike414, spike415, spike416, spike417, spike418, spike419, spike420, spike421, spike422, spike423, spike424, spike425, spike426, spike427, spike428, spike429, spike430, spike431, spike432, spike433, spike434, spike435, spike436, spike437, spike438, spike439, spike440, spike441, spike442, spike443, spike444, spike445, spike446, spike447, spike448, spike449) begin
        spike_register[400] = spike400;

        spike_register[401] = spike401;        spike_register[402] = spike402;        spike_register[403] = spike403;        spike_register[404] = spike404;        spike_register[405] = spike405;        spike_register[406] = spike406;        spike_register[407] = spike407;        spike_register[408] = spike408;        spike_register[409] = spike409;        spike_register[410] = spike410;        spike_register[411] = spike411;        spike_register[412] = spike412;        spike_register[413] = spike413;        spike_register[414] = spike414;        spike_register[415] = spike415;        spike_register[416] = spike416;        spike_register[417] = spike417;        spike_register[418] = spike418;        spike_register[419] = spike419;        spike_register[420] = spike420;        spike_register[421] = spike421;        spike_register[422] = spike422;        spike_register[423] = spike423;        spike_register[424] = spike424;        spike_register[425] = spike425;        spike_register[426] = spike426;        spike_register[427] = spike427;        spike_register[428] = spike428;        spike_register[429] = spike429;        spike_register[430] = spike430;        spike_register[431] = spike431;        spike_register[432] = spike432;        spike_register[433] = spike433;        spike_register[434] = spike434;        spike_register[435] = spike435;        spike_register[436] = spike436;        spike_register[437] = spike437;        spike_register[438] = spike438;        spike_register[439] = spike439;        spike_register[440] = spike440;        spike_register[441] = spike441;        spike_register[442] = spike442;        spike_register[443] = spike443;        spike_register[444] = spike444;        spike_register[445] = spike445;        spike_register[446] = spike446;        spike_register[447] = spike447;        spike_register[448] = spike448;        spike_register[449] = spike449;
        #0.5
        if(clear == 1'b0) begin
            for(i9 = 400; i9 <=449; i9= i9+1) begin
                if(spike_register[i9] == 1 && lock9 == 0) begin
                    lock9 = 1;
                    for(j9 = connection_pointer[i9]; j9 < connection_pointer[i9+1]; j9= j9+1) begin
                        packet9 = #0.1 {neuron_addresses[i9], downstream_connections[j9]};
                    end
                    spike_register[i9] = 0;
                    lock9 = 0;
                end
            end
        end

    end
    always @(clear, lock10, spike450, spike451, spike452, spike453, spike454, spike455, spike456, spike457, spike458, spike459, spike460, spike461, spike462, spike463, spike464, spike465, spike466, spike467, spike468, spike469, spike470, spike471, spike472, spike473, spike474, spike475, spike476, spike477, spike478, spike479, spike480, spike481, spike482, spike483, spike484, spike485, spike486, spike487, spike488, spike489, spike490, spike491, spike492, spike493, spike494, spike495, spike496, spike497, spike498, spike499) begin
        spike_register[450] = spike450;        spike_register[451] = spike451;        spike_register[452] = spike452;        spike_register[453] = spike453;        spike_register[454] = spike454;        spike_register[455] = spike455;        spike_register[456] = spike456;        spike_register[457] = spike457;        spike_register[458] = spike458;        spike_register[459] = spike459;        spike_register[460] = spike460;        spike_register[461] = spike461;        spike_register[462] = spike462;        spike_register[463] = spike463;        spike_register[464] = spike464;        spike_register[465] = spike465;        spike_register[466] = spike466;        spike_register[467] = spike467;        spike_register[468] = spike468;        spike_register[469] = spike469;        spike_register[470] = spike470;        spike_register[471] = spike471;        spike_register[472] = spike472;        spike_register[473] = spike473;        spike_register[474] = spike474;        spike_register[475] = spike475;        spike_register[476] = spike476;        spike_register[477] = spike477;        spike_register[478] = spike478;        spike_register[479] = spike479;        spike_register[480] = spike480;        spike_register[481] = spike481;        spike_register[482] = spike482;        spike_register[483] = spike483;        spike_register[484] = spike484;        spike_register[485] = spike485;        spike_register[486] = spike486;        spike_register[487] = spike487;        spike_register[488] = spike488;        spike_register[489] = spike489;        spike_register[490] = spike490;        spike_register[491] = spike491;        spike_register[492] = spike492;        spike_register[493] = spike493;        spike_register[494] = spike494;        spike_register[495] = spike495;        spike_register[496] = spike496;        spike_register[497] = spike497;        spike_register[498] = spike498;        spike_register[499] = spike499;
        #0.5
        if(clear == 1'b0) begin
            for(i10 = 450; i10 <=499; i10= i10+1) begin
                if(spike_register[i10] == 1 && lock10 == 0) begin
                    lock10 = 1;
                    for(j10 = connection_pointer[i10]; j10 < connection_pointer[i10+1]; j10= j10+1) begin
                        packet10 = #0.1 {neuron_addresses[i10], downstream_connections[j10]};
                    end
                    spike_register[i10] = 0;
                    lock10 = 0;
                end
            end
        end

    end
    always @(clear, lock11, spike500, spike501, spike502, spike503, spike504, spike505, spike506, spike507, spike508, spike509, spike510, spike511, spike512, spike513, spike514, spike515, spike516, spike517, spike518, spike519, spike520, spike521, spike522, spike523, spike524, spike525, spike526, spike527, spike528, spike529, spike530, spike531, spike532, spike533, spike534, spike535, spike536, spike537, spike538, spike539, spike540, spike541, spike542, spike543, spike544, spike545, spike546, spike547, spike548, spike549) begin
        spike_register[500] = spike500;

        spike_register[501] = spike501;        spike_register[502] = spike502;        spike_register[503] = spike503;        spike_register[504] = spike504;        spike_register[505] = spike505;        spike_register[506] = spike506;        spike_register[507] = spike507;        spike_register[508] = spike508;        spike_register[509] = spike509;        spike_register[510] = spike510;        spike_register[511] = spike511;        spike_register[512] = spike512;        spike_register[513] = spike513;        spike_register[514] = spike514;        spike_register[515] = spike515;        spike_register[516] = spike516;        spike_register[517] = spike517;        spike_register[518] = spike518;        spike_register[519] = spike519;        spike_register[520] = spike520;        spike_register[521] = spike521;        spike_register[522] = spike522;        spike_register[523] = spike523;        spike_register[524] = spike524;        spike_register[525] = spike525;        spike_register[526] = spike526;        spike_register[527] = spike527;        spike_register[528] = spike528;        spike_register[529] = spike529;        spike_register[530] = spike530;        spike_register[531] = spike531;        spike_register[532] = spike532;        spike_register[533] = spike533;        spike_register[534] = spike534;        spike_register[535] = spike535;        spike_register[536] = spike536;        spike_register[537] = spike537;        spike_register[538] = spike538;        spike_register[539] = spike539;        spike_register[540] = spike540;        spike_register[541] = spike541;        spike_register[542] = spike542;        spike_register[543] = spike543;        spike_register[544] = spike544;        spike_register[545] = spike545;        spike_register[546] = spike546;        spike_register[547] = spike547;        spike_register[548] = spike548;        spike_register[549] = spike549;
        #0.5
        if(clear == 1'b0) begin
            for(i11 = 500; i11 <=549; i11= i11+1) begin
                if(spike_register[i11] == 1 && lock11 == 0) begin
                    lock11 = 1;
                    for(j11 = connection_pointer[i11]; j11 < connection_pointer[i11+1]; j11= j11+1) begin
                        packet11 = #0.1 {neuron_addresses[i11], downstream_connections[j11]};
                    end
                    spike_register[i11] = 0;
                    lock11 = 0;
                end
            end
        end

    end
    always @(clear, lock12, spike550, spike551, spike552, spike553, spike554, spike555, spike556, spike557, spike558, spike559, spike560, spike561, spike562, spike563, spike564, spike565, spike566, spike567, spike568, spike569, spike570, spike571, spike572, spike573, spike574, spike575, spike576, spike577, spike578, spike579, spike580, spike581, spike582, spike583, spike584, spike585, spike586, spike587, spike588, spike589, spike590, spike591, spike592, spike593, spike594, spike595, spike596, spike597, spike598, spike599) begin
        spike_register[550] = spike550;        spike_register[551] = spike551;        spike_register[552] = spike552;        spike_register[553] = spike553;        spike_register[554] = spike554;        spike_register[555] = spike555;        spike_register[556] = spike556;        spike_register[557] = spike557;        spike_register[558] = spike558;        spike_register[559] = spike559;        spike_register[560] = spike560;        spike_register[561] = spike561;        spike_register[562] = spike562;        spike_register[563] = spike563;        spike_register[564] = spike564;        spike_register[565] = spike565;        spike_register[566] = spike566;        spike_register[567] = spike567;        spike_register[568] = spike568;        spike_register[569] = spike569;        spike_register[570] = spike570;        spike_register[571] = spike571;        spike_register[572] = spike572;        spike_register[573] = spike573;        spike_register[574] = spike574;        spike_register[575] = spike575;        spike_register[576] = spike576;        spike_register[577] = spike577;        spike_register[578] = spike578;        spike_register[579] = spike579;        spike_register[580] = spike580;        spike_register[581] = spike581;        spike_register[582] = spike582;        spike_register[583] = spike583;        spike_register[584] = spike584;        spike_register[585] = spike585;        spike_register[586] = spike586;        spike_register[587] = spike587;        spike_register[588] = spike588;        spike_register[589] = spike589;        spike_register[590] = spike590;        spike_register[591] = spike591;        spike_register[592] = spike592;        spike_register[593] = spike593;        spike_register[594] = spike594;        spike_register[595] = spike595;        spike_register[596] = spike596;        spike_register[597] = spike597;        spike_register[598] = spike598;        spike_register[599] = spike599;
        #0.5
        if(clear == 1'b0) begin
            for(i12 = 550; i12 <=599; i12= i12+1) begin
                if(spike_register[i12] == 1 && lock12 == 0) begin
                    lock12 = 1;
                    for(j12 = connection_pointer[i12]; j12 < connection_pointer[i12+1]; j12= j12+1) begin
                        packet12 = #0.1 {neuron_addresses[i12], downstream_connections[j12]};
                    end
                    spike_register[i12] = 0;
                    lock12 = 0;
                end
            end
        end

    end
    always @(clear, lock13, spike600, spike601, spike602, spike603, spike604, spike605, spike606, spike607, spike608, spike609, spike610, spike611, spike612, spike613, spike614, spike615, spike616, spike617, spike618, spike619, spike620, spike621, spike622, spike623, spike624, spike625, spike626, spike627, spike628, spike629, spike630, spike631, spike632, spike633, spike634, spike635, spike636, spike637, spike638, spike639, spike640, spike641, spike642, spike643, spike644, spike645, spike646, spike647, spike648, spike649) begin
        spike_register[600] = spike600;

        spike_register[601] = spike601;        spike_register[602] = spike602;        spike_register[603] = spike603;        spike_register[604] = spike604;        spike_register[605] = spike605;        spike_register[606] = spike606;        spike_register[607] = spike607;        spike_register[608] = spike608;        spike_register[609] = spike609;        spike_register[610] = spike610;        spike_register[611] = spike611;        spike_register[612] = spike612;        spike_register[613] = spike613;        spike_register[614] = spike614;        spike_register[615] = spike615;        spike_register[616] = spike616;        spike_register[617] = spike617;        spike_register[618] = spike618;        spike_register[619] = spike619;        spike_register[620] = spike620;        spike_register[621] = spike621;        spike_register[622] = spike622;        spike_register[623] = spike623;        spike_register[624] = spike624;        spike_register[625] = spike625;        spike_register[626] = spike626;        spike_register[627] = spike627;        spike_register[628] = spike628;        spike_register[629] = spike629;        spike_register[630] = spike630;        spike_register[631] = spike631;        spike_register[632] = spike632;        spike_register[633] = spike633;        spike_register[634] = spike634;        spike_register[635] = spike635;        spike_register[636] = spike636;        spike_register[637] = spike637;        spike_register[638] = spike638;        spike_register[639] = spike639;        spike_register[640] = spike640;        spike_register[641] = spike641;        spike_register[642] = spike642;        spike_register[643] = spike643;        spike_register[644] = spike644;        spike_register[645] = spike645;        spike_register[646] = spike646;        spike_register[647] = spike647;        spike_register[648] = spike648;        spike_register[649] = spike649;
        #0.5
        if(clear == 1'b0) begin
            for(i13 = 600; i13 <=649; i13= i13+1) begin
                if(spike_register[i13] == 1 && lock13 == 0) begin
                    lock13 = 1;
                    for(j13 = connection_pointer[i13]; j13 < connection_pointer[i13+1]; j13= j13+1) begin
                        packet13 = #0.1 {neuron_addresses[i13], downstream_connections[j13]};
                    end
                    spike_register[i13] = 0;
                    lock13 = 0;
                end
            end
        end

    end
    always @(clear, lock14, spike650, spike651, spike652, spike653, spike654, spike655, spike656, spike657, spike658, spike659, spike660, spike661, spike662, spike663, spike664, spike665, spike666, spike667, spike668, spike669, spike670, spike671, spike672, spike673, spike674, spike675, spike676, spike677, spike678, spike679, spike680, spike681, spike682, spike683, spike684, spike685, spike686, spike687, spike688, spike689, spike690, spike691, spike692, spike693, spike694, spike695, spike696, spike697, spike698, spike699) begin
        spike_register[650] = spike650;        spike_register[651] = spike651;        spike_register[652] = spike652;        spike_register[653] = spike653;        spike_register[654] = spike654;        spike_register[655] = spike655;        spike_register[656] = spike656;        spike_register[657] = spike657;        spike_register[658] = spike658;        spike_register[659] = spike659;        spike_register[660] = spike660;        spike_register[661] = spike661;        spike_register[662] = spike662;        spike_register[663] = spike663;        spike_register[664] = spike664;        spike_register[665] = spike665;        spike_register[666] = spike666;        spike_register[667] = spike667;        spike_register[668] = spike668;        spike_register[669] = spike669;        spike_register[670] = spike670;        spike_register[671] = spike671;        spike_register[672] = spike672;        spike_register[673] = spike673;        spike_register[674] = spike674;        spike_register[675] = spike675;        spike_register[676] = spike676;        spike_register[677] = spike677;        spike_register[678] = spike678;        spike_register[679] = spike679;        spike_register[680] = spike680;        spike_register[681] = spike681;        spike_register[682] = spike682;        spike_register[683] = spike683;        spike_register[684] = spike684;        spike_register[685] = spike685;        spike_register[686] = spike686;        spike_register[687] = spike687;        spike_register[688] = spike688;        spike_register[689] = spike689;        spike_register[690] = spike690;        spike_register[691] = spike691;        spike_register[692] = spike692;        spike_register[693] = spike693;        spike_register[694] = spike694;        spike_register[695] = spike695;        spike_register[696] = spike696;        spike_register[697] = spike697;        spike_register[698] = spike698;        spike_register[699] = spike699;
        #0.5
        if(clear == 1'b0) begin
            for(i14 = 650; i14 <=699; i14= i14+1) begin
                if(spike_register[i14] == 1 && lock14 == 0) begin
                    lock14 = 1;
                    for(j14 = connection_pointer[i14]; j14 < connection_pointer[i14+1]; j14= j14+1) begin
                        packet14 = #0.1 {neuron_addresses[i14], downstream_connections[j14]};
                    end
                    spike_register[i14] = 0;
                    lock14 = 0;
                end
            end
        end

    end
    always @(clear, lock15, spike700, spike701, spike702, spike703, spike704, spike705, spike706, spike707, spike708, spike709, spike710, spike711, spike712, spike713, spike714, spike715, spike716, spike717, spike718, spike719, spike720, spike721, spike722, spike723, spike724, spike725, spike726, spike727, spike728, spike729, spike730, spike731, spike732, spike733, spike734, spike735, spike736, spike737, spike738, spike739, spike740, spike741, spike742, spike743, spike744, spike745, spike746, spike747, spike748, spike749) begin
        spike_register[700] = spike700;

        spike_register[701] = spike701;        spike_register[702] = spike702;        spike_register[703] = spike703;        spike_register[704] = spike704;        spike_register[705] = spike705;        spike_register[706] = spike706;        spike_register[707] = spike707;        spike_register[708] = spike708;        spike_register[709] = spike709;        spike_register[710] = spike710;        spike_register[711] = spike711;        spike_register[712] = spike712;        spike_register[713] = spike713;        spike_register[714] = spike714;        spike_register[715] = spike715;        spike_register[716] = spike716;        spike_register[717] = spike717;        spike_register[718] = spike718;        spike_register[719] = spike719;        spike_register[720] = spike720;        spike_register[721] = spike721;        spike_register[722] = spike722;        spike_register[723] = spike723;        spike_register[724] = spike724;        spike_register[725] = spike725;        spike_register[726] = spike726;        spike_register[727] = spike727;        spike_register[728] = spike728;        spike_register[729] = spike729;        spike_register[730] = spike730;        spike_register[731] = spike731;        spike_register[732] = spike732;        spike_register[733] = spike733;        spike_register[734] = spike734;        spike_register[735] = spike735;        spike_register[736] = spike736;        spike_register[737] = spike737;        spike_register[738] = spike738;        spike_register[739] = spike739;        spike_register[740] = spike740;        spike_register[741] = spike741;        spike_register[742] = spike742;        spike_register[743] = spike743;        spike_register[744] = spike744;        spike_register[745] = spike745;        spike_register[746] = spike746;        spike_register[747] = spike747;        spike_register[748] = spike748;        spike_register[749] = spike749;
        #0.5
        if(clear == 1'b0) begin
            for(i15 = 700; i15 <=749; i15= i15+1) begin
                if(spike_register[i15] == 1 && lock15 == 0) begin
                    lock15 = 1;
                    for(j15 = connection_pointer[i15]; j15 < connection_pointer[i15+1]; j15= j15+1) begin
                        packet15 = #0.1 {neuron_addresses[i15], downstream_connections[j15]};
                    end
                    spike_register[i15] = 0;
                    lock15 = 0;
                end
            end
        end

    end
    always @(clear, lock16, spike750, spike751, spike752, spike753, spike754, spike755, spike756, spike757, spike758, spike759, spike760, spike761, spike762, spike763, spike764, spike765, spike766, spike767, spike768, spike769, spike770, spike771, spike772, spike773, spike774, spike775, spike776, spike777, spike778, spike779, spike780, spike781, spike782, spike783, spike784, spike785, spike786, spike787, spike788, spike789, spike790, spike791, spike792, spike793, spike794, spike795, spike796, spike797, spike798, spike799) begin
        spike_register[750] = spike750;        spike_register[751] = spike751;        spike_register[752] = spike752;        spike_register[753] = spike753;        spike_register[754] = spike754;        spike_register[755] = spike755;        spike_register[756] = spike756;        spike_register[757] = spike757;        spike_register[758] = spike758;        spike_register[759] = spike759;        spike_register[760] = spike760;        spike_register[761] = spike761;        spike_register[762] = spike762;        spike_register[763] = spike763;        spike_register[764] = spike764;        spike_register[765] = spike765;        spike_register[766] = spike766;        spike_register[767] = spike767;        spike_register[768] = spike768;        spike_register[769] = spike769;        spike_register[770] = spike770;        spike_register[771] = spike771;        spike_register[772] = spike772;        spike_register[773] = spike773;        spike_register[774] = spike774;        spike_register[775] = spike775;        spike_register[776] = spike776;        spike_register[777] = spike777;        spike_register[778] = spike778;        spike_register[779] = spike779;        spike_register[780] = spike780;        spike_register[781] = spike781;        spike_register[782] = spike782;        spike_register[783] = spike783;        spike_register[784] = spike784;        spike_register[785] = spike785;        spike_register[786] = spike786;        spike_register[787] = spike787;        spike_register[788] = spike788;        spike_register[789] = spike789;        spike_register[790] = spike790;        spike_register[791] = spike791;        spike_register[792] = spike792;        spike_register[793] = spike793;        spike_register[794] = spike794;        spike_register[795] = spike795;        spike_register[796] = spike796;        spike_register[797] = spike797;        spike_register[798] = spike798;        spike_register[799] = spike799;
        #0.5
        if(clear == 1'b0) begin
            for(i16 = 750; i16 <=799; i16= i16+1) begin
                if(spike_register[i16] == 1 && lock16 == 0) begin
                    lock16 = 1;
                    for(j16 = connection_pointer[i16]; j16 < connection_pointer[i16+1]; j16= j16+1) begin
                        packet16 = #0.1 {neuron_addresses[i16], downstream_connections[j16]};
                    end
                    spike_register[i16] = 0;
                    lock16 = 0;
                end
            end
        end

    end
    always @(clear, lock17, spike800, spike801, spike802, spike803, spike804, spike805, spike806, spike807, spike808, spike809, spike810, spike811, spike812, spike813, spike814, spike815, spike816, spike817, spike818, spike819, spike820, spike821, spike822, spike823, spike824, spike825, spike826, spike827, spike828, spike829, spike830, spike831, spike832, spike833, spike834, spike835, spike836, spike837, spike838, spike839, spike840, spike841, spike842, spike843, spike844, spike845, spike846, spike847, spike848, spike849) begin
        spike_register[800] = spike800;

        spike_register[801] = spike801;        spike_register[802] = spike802;        spike_register[803] = spike803;        spike_register[804] = spike804;        spike_register[805] = spike805;        spike_register[806] = spike806;        spike_register[807] = spike807;        spike_register[808] = spike808;        spike_register[809] = spike809;        spike_register[810] = spike810;        spike_register[811] = spike811;        spike_register[812] = spike812;        spike_register[813] = spike813;        spike_register[814] = spike814;        spike_register[815] = spike815;        spike_register[816] = spike816;        spike_register[817] = spike817;        spike_register[818] = spike818;        spike_register[819] = spike819;        spike_register[820] = spike820;        spike_register[821] = spike821;        spike_register[822] = spike822;        spike_register[823] = spike823;        spike_register[824] = spike824;        spike_register[825] = spike825;        spike_register[826] = spike826;        spike_register[827] = spike827;        spike_register[828] = spike828;        spike_register[829] = spike829;        spike_register[830] = spike830;        spike_register[831] = spike831;        spike_register[832] = spike832;        spike_register[833] = spike833;        spike_register[834] = spike834;        spike_register[835] = spike835;        spike_register[836] = spike836;        spike_register[837] = spike837;        spike_register[838] = spike838;        spike_register[839] = spike839;        spike_register[840] = spike840;        spike_register[841] = spike841;        spike_register[842] = spike842;        spike_register[843] = spike843;        spike_register[844] = spike844;        spike_register[845] = spike845;        spike_register[846] = spike846;        spike_register[847] = spike847;        spike_register[848] = spike848;        spike_register[849] = spike849;
        #0.5
        if(clear == 1'b0) begin
            for(i17 = 800; i17 <=849; i17= i17+1) begin
                if(spike_register[i17] == 1 && lock17 == 0) begin
                    lock17 = 1;
                    for(j17 = connection_pointer[i17]; j17 < connection_pointer[i17+1]; j17= j17+1) begin
                        packet17 = #0.1 {neuron_addresses[i17], downstream_connections[j17]};
                    end
                    spike_register[i17] = 0;
                    lock17 = 0;
                end
            end
        end

    end
    always @(clear, lock18, spike850, spike851, spike852, spike853, spike854, spike855, spike856, spike857, spike858, spike859, spike860, spike861, spike862, spike863, spike864, spike865, spike866, spike867, spike868, spike869, spike870, spike871, spike872, spike873, spike874, spike875, spike876, spike877, spike878, spike879, spike880, spike881, spike882, spike883, spike884, spike885, spike886, spike887, spike888, spike889, spike890, spike891, spike892, spike893, spike894, spike895, spike896, spike897, spike898, spike899) begin
        spike_register[850] = spike850;        spike_register[851] = spike851;        spike_register[852] = spike852;        spike_register[853] = spike853;        spike_register[854] = spike854;        spike_register[855] = spike855;        spike_register[856] = spike856;        spike_register[857] = spike857;        spike_register[858] = spike858;        spike_register[859] = spike859;        spike_register[860] = spike860;        spike_register[861] = spike861;        spike_register[862] = spike862;        spike_register[863] = spike863;        spike_register[864] = spike864;        spike_register[865] = spike865;        spike_register[866] = spike866;        spike_register[867] = spike867;        spike_register[868] = spike868;        spike_register[869] = spike869;        spike_register[870] = spike870;        spike_register[871] = spike871;        spike_register[872] = spike872;        spike_register[873] = spike873;        spike_register[874] = spike874;        spike_register[875] = spike875;        spike_register[876] = spike876;        spike_register[877] = spike877;        spike_register[878] = spike878;        spike_register[879] = spike879;        spike_register[880] = spike880;        spike_register[881] = spike881;        spike_register[882] = spike882;        spike_register[883] = spike883;        spike_register[884] = spike884;        spike_register[885] = spike885;        spike_register[886] = spike886;        spike_register[887] = spike887;        spike_register[888] = spike888;        spike_register[889] = spike889;        spike_register[890] = spike890;        spike_register[891] = spike891;        spike_register[892] = spike892;        spike_register[893] = spike893;        spike_register[894] = spike894;        spike_register[895] = spike895;        spike_register[896] = spike896;        spike_register[897] = spike897;        spike_register[898] = spike898;        spike_register[899] = spike899;
        #0.5
        if(clear == 1'b0) begin
            for(i18 = 850; i18 <=899; i18= i18+1) begin
                if(spike_register[i18] == 1 && lock18 == 0) begin
                    lock18 = 1;
                    for(j18 = connection_pointer[i18]; j18 < connection_pointer[i18+1]; j18= j18+1) begin
                        packet18 = #0.1 {neuron_addresses[i18], downstream_connections[j18]};
                    end
                    spike_register[i18] = 0;
                    lock18 = 0;
                end
            end
        end

    end
    always @(clear, lock19, spike900, spike901, spike902, spike903, spike904, spike905, spike906, spike907, spike908, spike909, spike910, spike911, spike912, spike913, spike914, spike915, spike916, spike917, spike918, spike919, spike920, spike921, spike922, spike923, spike924, spike925, spike926, spike927, spike928, spike929, spike930, spike931, spike932, spike933, spike934, spike935, spike936, spike937, spike938, spike939, spike940, spike941, spike942, spike943, spike944, spike945, spike946, spike947, spike948, spike949) begin
        spike_register[900] = spike900;

        spike_register[901] = spike901;        spike_register[902] = spike902;        spike_register[903] = spike903;        spike_register[904] = spike904;        spike_register[905] = spike905;        spike_register[906] = spike906;        spike_register[907] = spike907;        spike_register[908] = spike908;        spike_register[909] = spike909;        spike_register[910] = spike910;        spike_register[911] = spike911;        spike_register[912] = spike912;        spike_register[913] = spike913;        spike_register[914] = spike914;        spike_register[915] = spike915;        spike_register[916] = spike916;        spike_register[917] = spike917;        spike_register[918] = spike918;        spike_register[919] = spike919;        spike_register[920] = spike920;        spike_register[921] = spike921;        spike_register[922] = spike922;        spike_register[923] = spike923;        spike_register[924] = spike924;        spike_register[925] = spike925;        spike_register[926] = spike926;        spike_register[927] = spike927;        spike_register[928] = spike928;        spike_register[929] = spike929;        spike_register[930] = spike930;        spike_register[931] = spike931;        spike_register[932] = spike932;        spike_register[933] = spike933;        spike_register[934] = spike934;        spike_register[935] = spike935;        spike_register[936] = spike936;        spike_register[937] = spike937;        spike_register[938] = spike938;        spike_register[939] = spike939;        spike_register[940] = spike940;        spike_register[941] = spike941;        spike_register[942] = spike942;        spike_register[943] = spike943;        spike_register[944] = spike944;        spike_register[945] = spike945;        spike_register[946] = spike946;        spike_register[947] = spike947;        spike_register[948] = spike948;        spike_register[949] = spike949;
        #0.5
        if(clear == 1'b0) begin
            for(i19 = 900; i19 <=949; i19= i19+1) begin
                if(spike_register[i19] == 1 && lock19 == 0) begin
                    lock19 = 1;
                    for(j19 = connection_pointer[i19]; j19 < connection_pointer[i19+1]; j19= j19+1) begin
                        packet19 = #0.1 {neuron_addresses[i19], downstream_connections[j19]};
                    end
                    spike_register[i19] = 0;
                    lock19 = 0;
                end
            end
        end

    end
    always @(clear, lock20, spike950, spike951, spike952, spike953, spike954, spike955, spike956, spike957, spike958, spike959, spike960, spike961, spike962, spike963, spike964, spike965, spike966, spike967, spike968, spike969, spike970, spike971, spike972, spike973, spike974, spike975, spike976, spike977, spike978, spike979, spike980, spike981, spike982, spike983, spike984, spike985, spike986, spike987, spike988, spike989, spike990, spike991, spike992, spike993, spike994, spike995, spike996, spike997, spike998, spike999) begin
        spike_register[950] = spike950;        spike_register[951] = spike951;        spike_register[952] = spike952;        spike_register[953] = spike953;        spike_register[954] = spike954;        spike_register[955] = spike955;        spike_register[956] = spike956;        spike_register[957] = spike957;        spike_register[958] = spike958;        spike_register[959] = spike959;        spike_register[960] = spike960;        spike_register[961] = spike961;        spike_register[962] = spike962;        spike_register[963] = spike963;        spike_register[964] = spike964;        spike_register[965] = spike965;        spike_register[966] = spike966;        spike_register[967] = spike967;        spike_register[968] = spike968;        spike_register[969] = spike969;        spike_register[970] = spike970;        spike_register[971] = spike971;        spike_register[972] = spike972;        spike_register[973] = spike973;        spike_register[974] = spike974;        spike_register[975] = spike975;        spike_register[976] = spike976;        spike_register[977] = spike977;        spike_register[978] = spike978;        spike_register[979] = spike979;        spike_register[980] = spike980;        spike_register[981] = spike981;        spike_register[982] = spike982;        spike_register[983] = spike983;        spike_register[984] = spike984;        spike_register[985] = spike985;        spike_register[986] = spike986;        spike_register[987] = spike987;        spike_register[988] = spike988;        spike_register[989] = spike989;        spike_register[990] = spike990;        spike_register[991] = spike991;        spike_register[992] = spike992;        spike_register[993] = spike993;        spike_register[994] = spike994;        spike_register[995] = spike995;        spike_register[996] = spike996;        spike_register[997] = spike997;        spike_register[998] = spike998;        spike_register[999] = spike999;
        #0.5
        if(clear == 1'b0) begin
            for(i20 = 950; i20 <=999; i20= i20+1) begin
                if(spike_register[i20] == 1 && lock20 == 0) begin
                    lock20 = 1;
                    for(j20 = connection_pointer[i20]; j20 < connection_pointer[i20+1]; j20= j20+1) begin
                        packet20 = #0.1 {neuron_addresses[i20], downstream_connections[j20]};
                    end
                    spike_register[i20] = 0;
                    lock20 = 0;
                end
            end
        end

    end
    always @(clear, lock21, spike1000, spike1001, spike1002, spike1003, spike1004, spike1005, spike1006, spike1007, spike1008, spike1009, spike1010, spike1011, spike1012, spike1013, spike1014, spike1015, spike1016, spike1017, spike1018, spike1019, spike1020, spike1021, spike1022, spike1023) begin
        spike_register[1000] = spike1000;

        spike_register[1001] = spike1001;        spike_register[1002] = spike1002;        spike_register[1003] = spike1003;        spike_register[1004] = spike1004;        spike_register[1005] = spike1005;        spike_register[1006] = spike1006;        spike_register[1007] = spike1007;        spike_register[1008] = spike1008;        spike_register[1009] = spike1009;        spike_register[1010] = spike1010;        spike_register[1011] = spike1011;        spike_register[1012] = spike1012;        spike_register[1013] = spike1013;        spike_register[1014] = spike1014;        spike_register[1015] = spike1015;        spike_register[1016] = spike1016;        spike_register[1017] = spike1017;        spike_register[1018] = spike1018;        spike_register[1019] = spike1019;        spike_register[1020] = spike1020;        spike_register[1021] = spike1021;        spike_register[1022] = spike1022;        spike_register[1023] = spike1023;
        #0.5
        if(clear == 1'b0) begin
            for(i21 = 1000; i21 <=1049; i21= i21+1) begin
                if(spike_register[i21] == 1 && lock21 == 0) begin
                    lock21 = 1;
                    for(j21 = connection_pointer[i21]; j21 < connection_pointer[i21+1]; j21= j21+1) begin
                        packet21 = #0.1 {neuron_addresses[i21], downstream_connections[j21]};
                    end
                    spike_register[i21] = 0;
                    lock21 = 0;
                end
            end
        end

    end
    always @(packet1) begin 
        spike_origin = packet1[23:12];
        spike_destination = packet1[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet2) begin 
        spike_origin = packet2[23:12];
        spike_destination = packet2[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet3) begin 
        spike_origin = packet3[23:12];
        spike_destination = packet3[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet4) begin 
        spike_origin = packet4[23:12];
        spike_destination = packet4[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet5) begin 
        spike_origin = packet5[23:12];
        spike_destination = packet5[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet6) begin 
        spike_origin = packet6[23:12];
        spike_destination = packet6[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet7) begin 
        spike_origin = packet7[23:12];
        spike_destination = packet7[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet8) begin 
        spike_origin = packet8[23:12];
        spike_destination = packet8[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet9) begin 
        spike_origin = packet9[23:12];
        spike_destination = packet9[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet10) begin 
        spike_origin = packet10[23:12];
        spike_destination = packet10[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet11) begin 
        spike_origin = packet11[23:12];
        spike_destination = packet11[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet12) begin 
        spike_origin = packet12[23:12];
        spike_destination = packet12[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet13) begin 
        spike_origin = packet13[23:12];
        spike_destination = packet13[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet14) begin 
        spike_origin = packet14[23:12];
        spike_destination = packet14[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet15) begin 
        spike_origin = packet15[23:12];
        spike_destination = packet15[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet16) begin 
        spike_origin = packet16[23:12];
        spike_destination = packet16[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet17) begin 
        spike_origin = packet17[23:12];
        spike_destination = packet17[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet18) begin 
        spike_origin = packet18[23:12];
        spike_destination = packet18[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet19) begin 
        spike_origin = packet19[23:12];
        spike_destination = packet19[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet20) begin 
        spike_origin = packet20[23:12];
        spike_destination = packet20[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet21) begin 
        spike_origin = packet21[23:12];
        spike_destination = packet21[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(spike_out_source_array[0]) begin 
        spike_out_source0 = spike_out_source_array[0];
    end
    always @(spike_out_source_array[1]) begin 
        spike_out_source1 = spike_out_source_array[1];
    end
    always @(spike_out_source_array[2]) begin 
        spike_out_source2 = spike_out_source_array[2];
    end
    always @(spike_out_source_array[3]) begin 
        spike_out_source3 = spike_out_source_array[3];
    end
    always @(spike_out_source_array[4]) begin 
        spike_out_source4 = spike_out_source_array[4];
    end
    always @(spike_out_source_array[5]) begin 
        spike_out_source5 = spike_out_source_array[5];
    end
    always @(spike_out_source_array[6]) begin 
        spike_out_source6 = spike_out_source_array[6];
    end
    always @(spike_out_source_array[7]) begin 
        spike_out_source7 = spike_out_source_array[7];
    end
    always @(spike_out_source_array[8]) begin 
        spike_out_source8 = spike_out_source_array[8];
    end
    always @(spike_out_source_array[9]) begin 
        spike_out_source9 = spike_out_source_array[9];
    end
    always @(spike_out_source_array[10]) begin 
        spike_out_source10 = spike_out_source_array[10];
    end
    always @(spike_out_source_array[11]) begin 
        spike_out_source11 = spike_out_source_array[11];
    end
    always @(spike_out_source_array[12]) begin 
        spike_out_source12 = spike_out_source_array[12];
    end
    always @(spike_out_source_array[13]) begin 
        spike_out_source13 = spike_out_source_array[13];
    end
    always @(spike_out_source_array[14]) begin 
        spike_out_source14 = spike_out_source_array[14];
    end
    always @(spike_out_source_array[15]) begin 
        spike_out_source15 = spike_out_source_array[15];
    end
    always @(spike_out_source_array[16]) begin 
        spike_out_source16 = spike_out_source_array[16];
    end
    always @(spike_out_source_array[17]) begin 
        spike_out_source17 = spike_out_source_array[17];
    end
    always @(spike_out_source_array[18]) begin 
        spike_out_source18 = spike_out_source_array[18];
    end
    always @(spike_out_source_array[19]) begin 
        spike_out_source19 = spike_out_source_array[19];
    end
    always @(spike_out_source_array[20]) begin 
        spike_out_source20 = spike_out_source_array[20];
    end
    always @(spike_out_source_array[21]) begin 
        spike_out_source21 = spike_out_source_array[21];
    end
    always @(spike_out_source_array[22]) begin 
        spike_out_source22 = spike_out_source_array[22];
    end
    always @(spike_out_source_array[23]) begin 
        spike_out_source23 = spike_out_source_array[23];
    end
    always @(spike_out_source_array[24]) begin 
        spike_out_source24 = spike_out_source_array[24];
    end
    always @(spike_out_source_array[25]) begin 
        spike_out_source25 = spike_out_source_array[25];
    end
    always @(spike_out_source_array[26]) begin 
        spike_out_source26 = spike_out_source_array[26];
    end
    always @(spike_out_source_array[27]) begin 
        spike_out_source27 = spike_out_source_array[27];
    end
    always @(spike_out_source_array[28]) begin 
        spike_out_source28 = spike_out_source_array[28];
    end
    always @(spike_out_source_array[29]) begin 
        spike_out_source29 = spike_out_source_array[29];
    end
    always @(spike_out_source_array[30]) begin 
        spike_out_source30 = spike_out_source_array[30];
    end
    always @(spike_out_source_array[31]) begin 
        spike_out_source31 = spike_out_source_array[31];
    end
    always @(spike_out_source_array[32]) begin 
        spike_out_source32 = spike_out_source_array[32];
    end
    always @(spike_out_source_array[33]) begin 
        spike_out_source33 = spike_out_source_array[33];
    end
    always @(spike_out_source_array[34]) begin 
        spike_out_source34 = spike_out_source_array[34];
    end
    always @(spike_out_source_array[35]) begin 
        spike_out_source35 = spike_out_source_array[35];
    end
    always @(spike_out_source_array[36]) begin 
        spike_out_source36 = spike_out_source_array[36];
    end
    always @(spike_out_source_array[37]) begin 
        spike_out_source37 = spike_out_source_array[37];
    end
    always @(spike_out_source_array[38]) begin 
        spike_out_source38 = spike_out_source_array[38];
    end
    always @(spike_out_source_array[39]) begin 
        spike_out_source39 = spike_out_source_array[39];
    end
    always @(spike_out_source_array[40]) begin 
        spike_out_source40 = spike_out_source_array[40];
    end
    always @(spike_out_source_array[41]) begin 
        spike_out_source41 = spike_out_source_array[41];
    end
    always @(spike_out_source_array[42]) begin 
        spike_out_source42 = spike_out_source_array[42];
    end
    always @(spike_out_source_array[43]) begin 
        spike_out_source43 = spike_out_source_array[43];
    end
    always @(spike_out_source_array[44]) begin 
        spike_out_source44 = spike_out_source_array[44];
    end
    always @(spike_out_source_array[45]) begin 
        spike_out_source45 = spike_out_source_array[45];
    end
    always @(spike_out_source_array[46]) begin 
        spike_out_source46 = spike_out_source_array[46];
    end
    always @(spike_out_source_array[47]) begin 
        spike_out_source47 = spike_out_source_array[47];
    end
    always @(spike_out_source_array[48]) begin 
        spike_out_source48 = spike_out_source_array[48];
    end
    always @(spike_out_source_array[49]) begin 
        spike_out_source49 = spike_out_source_array[49];
    end
    always @(spike_out_source_array[50]) begin 
        spike_out_source50 = spike_out_source_array[50];
    end
    always @(spike_out_source_array[51]) begin 
        spike_out_source51 = spike_out_source_array[51];
    end
    always @(spike_out_source_array[52]) begin 
        spike_out_source52 = spike_out_source_array[52];
    end
    always @(spike_out_source_array[53]) begin 
        spike_out_source53 = spike_out_source_array[53];
    end
    always @(spike_out_source_array[54]) begin 
        spike_out_source54 = spike_out_source_array[54];
    end
    always @(spike_out_source_array[55]) begin 
        spike_out_source55 = spike_out_source_array[55];
    end
    always @(spike_out_source_array[56]) begin 
        spike_out_source56 = spike_out_source_array[56];
    end
    always @(spike_out_source_array[57]) begin 
        spike_out_source57 = spike_out_source_array[57];
    end
    always @(spike_out_source_array[58]) begin 
        spike_out_source58 = spike_out_source_array[58];
    end
    always @(spike_out_source_array[59]) begin 
        spike_out_source59 = spike_out_source_array[59];
    end
    always @(spike_out_source_array[60]) begin 
        spike_out_source60 = spike_out_source_array[60];
    end
    always @(spike_out_source_array[61]) begin 
        spike_out_source61 = spike_out_source_array[61];
    end
    always @(spike_out_source_array[62]) begin 
        spike_out_source62 = spike_out_source_array[62];
    end
    always @(spike_out_source_array[63]) begin 
        spike_out_source63 = spike_out_source_array[63];
    end
    always @(spike_out_source_array[64]) begin 
        spike_out_source64 = spike_out_source_array[64];
    end
    always @(spike_out_source_array[65]) begin 
        spike_out_source65 = spike_out_source_array[65];
    end
    always @(spike_out_source_array[66]) begin 
        spike_out_source66 = spike_out_source_array[66];
    end
    always @(spike_out_source_array[67]) begin 
        spike_out_source67 = spike_out_source_array[67];
    end
    always @(spike_out_source_array[68]) begin 
        spike_out_source68 = spike_out_source_array[68];
    end
    always @(spike_out_source_array[69]) begin 
        spike_out_source69 = spike_out_source_array[69];
    end
    always @(spike_out_source_array[70]) begin 
        spike_out_source70 = spike_out_source_array[70];
    end
    always @(spike_out_source_array[71]) begin 
        spike_out_source71 = spike_out_source_array[71];
    end
    always @(spike_out_source_array[72]) begin 
        spike_out_source72 = spike_out_source_array[72];
    end
    always @(spike_out_source_array[73]) begin 
        spike_out_source73 = spike_out_source_array[73];
    end
    always @(spike_out_source_array[74]) begin 
        spike_out_source74 = spike_out_source_array[74];
    end
    always @(spike_out_source_array[75]) begin 
        spike_out_source75 = spike_out_source_array[75];
    end
    always @(spike_out_source_array[76]) begin 
        spike_out_source76 = spike_out_source_array[76];
    end
    always @(spike_out_source_array[77]) begin 
        spike_out_source77 = spike_out_source_array[77];
    end
    always @(spike_out_source_array[78]) begin 
        spike_out_source78 = spike_out_source_array[78];
    end
    always @(spike_out_source_array[79]) begin 
        spike_out_source79 = spike_out_source_array[79];
    end
    always @(spike_out_source_array[80]) begin 
        spike_out_source80 = spike_out_source_array[80];
    end
    always @(spike_out_source_array[81]) begin 
        spike_out_source81 = spike_out_source_array[81];
    end
    always @(spike_out_source_array[82]) begin 
        spike_out_source82 = spike_out_source_array[82];
    end
    always @(spike_out_source_array[83]) begin 
        spike_out_source83 = spike_out_source_array[83];
    end
    always @(spike_out_source_array[84]) begin 
        spike_out_source84 = spike_out_source_array[84];
    end
    always @(spike_out_source_array[85]) begin 
        spike_out_source85 = spike_out_source_array[85];
    end
    always @(spike_out_source_array[86]) begin 
        spike_out_source86 = spike_out_source_array[86];
    end
    always @(spike_out_source_array[87]) begin 
        spike_out_source87 = spike_out_source_array[87];
    end
    always @(spike_out_source_array[88]) begin 
        spike_out_source88 = spike_out_source_array[88];
    end
    always @(spike_out_source_array[89]) begin 
        spike_out_source89 = spike_out_source_array[89];
    end
    always @(spike_out_source_array[90]) begin 
        spike_out_source90 = spike_out_source_array[90];
    end
    always @(spike_out_source_array[91]) begin 
        spike_out_source91 = spike_out_source_array[91];
    end
    always @(spike_out_source_array[92]) begin 
        spike_out_source92 = spike_out_source_array[92];
    end
    always @(spike_out_source_array[93]) begin 
        spike_out_source93 = spike_out_source_array[93];
    end
    always @(spike_out_source_array[94]) begin 
        spike_out_source94 = spike_out_source_array[94];
    end
    always @(spike_out_source_array[95]) begin 
        spike_out_source95 = spike_out_source_array[95];
    end
    always @(spike_out_source_array[96]) begin 
        spike_out_source96 = spike_out_source_array[96];
    end
    always @(spike_out_source_array[97]) begin 
        spike_out_source97 = spike_out_source_array[97];
    end
    always @(spike_out_source_array[98]) begin 
        spike_out_source98 = spike_out_source_array[98];
    end
    always @(spike_out_source_array[99]) begin 
        spike_out_source99 = spike_out_source_array[99];
    end
    always @(spike_out_source_array[100]) begin 
        spike_out_source100 = spike_out_source_array[100];
    end
    always @(spike_out_source_array[101]) begin 
        spike_out_source101 = spike_out_source_array[101];
    end
    always @(spike_out_source_array[102]) begin 
        spike_out_source102 = spike_out_source_array[102];
    end
    always @(spike_out_source_array[103]) begin 
        spike_out_source103 = spike_out_source_array[103];
    end
    always @(spike_out_source_array[104]) begin 
        spike_out_source104 = spike_out_source_array[104];
    end
    always @(spike_out_source_array[105]) begin 
        spike_out_source105 = spike_out_source_array[105];
    end
    always @(spike_out_source_array[106]) begin 
        spike_out_source106 = spike_out_source_array[106];
    end
    always @(spike_out_source_array[107]) begin 
        spike_out_source107 = spike_out_source_array[107];
    end
    always @(spike_out_source_array[108]) begin 
        spike_out_source108 = spike_out_source_array[108];
    end
    always @(spike_out_source_array[109]) begin 
        spike_out_source109 = spike_out_source_array[109];
    end
    always @(spike_out_source_array[110]) begin 
        spike_out_source110 = spike_out_source_array[110];
    end
    always @(spike_out_source_array[111]) begin 
        spike_out_source111 = spike_out_source_array[111];
    end
    always @(spike_out_source_array[112]) begin 
        spike_out_source112 = spike_out_source_array[112];
    end
    always @(spike_out_source_array[113]) begin 
        spike_out_source113 = spike_out_source_array[113];
    end
    always @(spike_out_source_array[114]) begin 
        spike_out_source114 = spike_out_source_array[114];
    end
    always @(spike_out_source_array[115]) begin 
        spike_out_source115 = spike_out_source_array[115];
    end
    always @(spike_out_source_array[116]) begin 
        spike_out_source116 = spike_out_source_array[116];
    end
    always @(spike_out_source_array[117]) begin 
        spike_out_source117 = spike_out_source_array[117];
    end
    always @(spike_out_source_array[118]) begin 
        spike_out_source118 = spike_out_source_array[118];
    end
    always @(spike_out_source_array[119]) begin 
        spike_out_source119 = spike_out_source_array[119];
    end
    always @(spike_out_source_array[120]) begin 
        spike_out_source120 = spike_out_source_array[120];
    end
    always @(spike_out_source_array[121]) begin 
        spike_out_source121 = spike_out_source_array[121];
    end
    always @(spike_out_source_array[122]) begin 
        spike_out_source122 = spike_out_source_array[122];
    end
    always @(spike_out_source_array[123]) begin 
        spike_out_source123 = spike_out_source_array[123];
    end
    always @(spike_out_source_array[124]) begin 
        spike_out_source124 = spike_out_source_array[124];
    end
    always @(spike_out_source_array[125]) begin 
        spike_out_source125 = spike_out_source_array[125];
    end
    always @(spike_out_source_array[126]) begin 
        spike_out_source126 = spike_out_source_array[126];
    end
    always @(spike_out_source_array[127]) begin 
        spike_out_source127 = spike_out_source_array[127];
    end
    always @(spike_out_source_array[128]) begin 
        spike_out_source128 = spike_out_source_array[128];
    end
    always @(spike_out_source_array[129]) begin 
        spike_out_source129 = spike_out_source_array[129];
    end
    always @(spike_out_source_array[130]) begin 
        spike_out_source130 = spike_out_source_array[130];
    end
    always @(spike_out_source_array[131]) begin 
        spike_out_source131 = spike_out_source_array[131];
    end
    always @(spike_out_source_array[132]) begin 
        spike_out_source132 = spike_out_source_array[132];
    end
    always @(spike_out_source_array[133]) begin 
        spike_out_source133 = spike_out_source_array[133];
    end
    always @(spike_out_source_array[134]) begin 
        spike_out_source134 = spike_out_source_array[134];
    end
    always @(spike_out_source_array[135]) begin 
        spike_out_source135 = spike_out_source_array[135];
    end
    always @(spike_out_source_array[136]) begin 
        spike_out_source136 = spike_out_source_array[136];
    end
    always @(spike_out_source_array[137]) begin 
        spike_out_source137 = spike_out_source_array[137];
    end
    always @(spike_out_source_array[138]) begin 
        spike_out_source138 = spike_out_source_array[138];
    end
    always @(spike_out_source_array[139]) begin 
        spike_out_source139 = spike_out_source_array[139];
    end
    always @(spike_out_source_array[140]) begin 
        spike_out_source140 = spike_out_source_array[140];
    end
    always @(spike_out_source_array[141]) begin 
        spike_out_source141 = spike_out_source_array[141];
    end
    always @(spike_out_source_array[142]) begin 
        spike_out_source142 = spike_out_source_array[142];
    end
    always @(spike_out_source_array[143]) begin 
        spike_out_source143 = spike_out_source_array[143];
    end
    always @(spike_out_source_array[144]) begin 
        spike_out_source144 = spike_out_source_array[144];
    end
    always @(spike_out_source_array[145]) begin 
        spike_out_source145 = spike_out_source_array[145];
    end
    always @(spike_out_source_array[146]) begin 
        spike_out_source146 = spike_out_source_array[146];
    end
    always @(spike_out_source_array[147]) begin 
        spike_out_source147 = spike_out_source_array[147];
    end
    always @(spike_out_source_array[148]) begin 
        spike_out_source148 = spike_out_source_array[148];
    end
    always @(spike_out_source_array[149]) begin 
        spike_out_source149 = spike_out_source_array[149];
    end
    always @(spike_out_source_array[150]) begin 
        spike_out_source150 = spike_out_source_array[150];
    end
    always @(spike_out_source_array[151]) begin 
        spike_out_source151 = spike_out_source_array[151];
    end
    always @(spike_out_source_array[152]) begin 
        spike_out_source152 = spike_out_source_array[152];
    end
    always @(spike_out_source_array[153]) begin 
        spike_out_source153 = spike_out_source_array[153];
    end
    always @(spike_out_source_array[154]) begin 
        spike_out_source154 = spike_out_source_array[154];
    end
    always @(spike_out_source_array[155]) begin 
        spike_out_source155 = spike_out_source_array[155];
    end
    always @(spike_out_source_array[156]) begin 
        spike_out_source156 = spike_out_source_array[156];
    end
    always @(spike_out_source_array[157]) begin 
        spike_out_source157 = spike_out_source_array[157];
    end
    always @(spike_out_source_array[158]) begin 
        spike_out_source158 = spike_out_source_array[158];
    end
    always @(spike_out_source_array[159]) begin 
        spike_out_source159 = spike_out_source_array[159];
    end
    always @(spike_out_source_array[160]) begin 
        spike_out_source160 = spike_out_source_array[160];
    end
    always @(spike_out_source_array[161]) begin 
        spike_out_source161 = spike_out_source_array[161];
    end
    always @(spike_out_source_array[162]) begin 
        spike_out_source162 = spike_out_source_array[162];
    end
    always @(spike_out_source_array[163]) begin 
        spike_out_source163 = spike_out_source_array[163];
    end
    always @(spike_out_source_array[164]) begin 
        spike_out_source164 = spike_out_source_array[164];
    end
    always @(spike_out_source_array[165]) begin 
        spike_out_source165 = spike_out_source_array[165];
    end
    always @(spike_out_source_array[166]) begin 
        spike_out_source166 = spike_out_source_array[166];
    end
    always @(spike_out_source_array[167]) begin 
        spike_out_source167 = spike_out_source_array[167];
    end
    always @(spike_out_source_array[168]) begin 
        spike_out_source168 = spike_out_source_array[168];
    end
    always @(spike_out_source_array[169]) begin 
        spike_out_source169 = spike_out_source_array[169];
    end
    always @(spike_out_source_array[170]) begin 
        spike_out_source170 = spike_out_source_array[170];
    end
    always @(spike_out_source_array[171]) begin 
        spike_out_source171 = spike_out_source_array[171];
    end
    always @(spike_out_source_array[172]) begin 
        spike_out_source172 = spike_out_source_array[172];
    end
    always @(spike_out_source_array[173]) begin 
        spike_out_source173 = spike_out_source_array[173];
    end
    always @(spike_out_source_array[174]) begin 
        spike_out_source174 = spike_out_source_array[174];
    end
    always @(spike_out_source_array[175]) begin 
        spike_out_source175 = spike_out_source_array[175];
    end
    always @(spike_out_source_array[176]) begin 
        spike_out_source176 = spike_out_source_array[176];
    end
    always @(spike_out_source_array[177]) begin 
        spike_out_source177 = spike_out_source_array[177];
    end
    always @(spike_out_source_array[178]) begin 
        spike_out_source178 = spike_out_source_array[178];
    end
    always @(spike_out_source_array[179]) begin 
        spike_out_source179 = spike_out_source_array[179];
    end
    always @(spike_out_source_array[180]) begin 
        spike_out_source180 = spike_out_source_array[180];
    end
    always @(spike_out_source_array[181]) begin 
        spike_out_source181 = spike_out_source_array[181];
    end
    always @(spike_out_source_array[182]) begin 
        spike_out_source182 = spike_out_source_array[182];
    end
    always @(spike_out_source_array[183]) begin 
        spike_out_source183 = spike_out_source_array[183];
    end
    always @(spike_out_source_array[184]) begin 
        spike_out_source184 = spike_out_source_array[184];
    end
    always @(spike_out_source_array[185]) begin 
        spike_out_source185 = spike_out_source_array[185];
    end
    always @(spike_out_source_array[186]) begin 
        spike_out_source186 = spike_out_source_array[186];
    end
    always @(spike_out_source_array[187]) begin 
        spike_out_source187 = spike_out_source_array[187];
    end
    always @(spike_out_source_array[188]) begin 
        spike_out_source188 = spike_out_source_array[188];
    end
    always @(spike_out_source_array[189]) begin 
        spike_out_source189 = spike_out_source_array[189];
    end
    always @(spike_out_source_array[190]) begin 
        spike_out_source190 = spike_out_source_array[190];
    end
    always @(spike_out_source_array[191]) begin 
        spike_out_source191 = spike_out_source_array[191];
    end
    always @(spike_out_source_array[192]) begin 
        spike_out_source192 = spike_out_source_array[192];
    end
    always @(spike_out_source_array[193]) begin 
        spike_out_source193 = spike_out_source_array[193];
    end
    always @(spike_out_source_array[194]) begin 
        spike_out_source194 = spike_out_source_array[194];
    end
    always @(spike_out_source_array[195]) begin 
        spike_out_source195 = spike_out_source_array[195];
    end
    always @(spike_out_source_array[196]) begin 
        spike_out_source196 = spike_out_source_array[196];
    end
    always @(spike_out_source_array[197]) begin 
        spike_out_source197 = spike_out_source_array[197];
    end
    always @(spike_out_source_array[198]) begin 
        spike_out_source198 = spike_out_source_array[198];
    end
    always @(spike_out_source_array[199]) begin 
        spike_out_source199 = spike_out_source_array[199];
    end
    always @(spike_out_source_array[200]) begin 
        spike_out_source200 = spike_out_source_array[200];
    end
    always @(spike_out_source_array[201]) begin 
        spike_out_source201 = spike_out_source_array[201];
    end
    always @(spike_out_source_array[202]) begin 
        spike_out_source202 = spike_out_source_array[202];
    end
    always @(spike_out_source_array[203]) begin 
        spike_out_source203 = spike_out_source_array[203];
    end
    always @(spike_out_source_array[204]) begin 
        spike_out_source204 = spike_out_source_array[204];
    end
    always @(spike_out_source_array[205]) begin 
        spike_out_source205 = spike_out_source_array[205];
    end
    always @(spike_out_source_array[206]) begin 
        spike_out_source206 = spike_out_source_array[206];
    end
    always @(spike_out_source_array[207]) begin 
        spike_out_source207 = spike_out_source_array[207];
    end
    always @(spike_out_source_array[208]) begin 
        spike_out_source208 = spike_out_source_array[208];
    end
    always @(spike_out_source_array[209]) begin 
        spike_out_source209 = spike_out_source_array[209];
    end
    always @(spike_out_source_array[210]) begin 
        spike_out_source210 = spike_out_source_array[210];
    end
    always @(spike_out_source_array[211]) begin 
        spike_out_source211 = spike_out_source_array[211];
    end
    always @(spike_out_source_array[212]) begin 
        spike_out_source212 = spike_out_source_array[212];
    end
    always @(spike_out_source_array[213]) begin 
        spike_out_source213 = spike_out_source_array[213];
    end
    always @(spike_out_source_array[214]) begin 
        spike_out_source214 = spike_out_source_array[214];
    end
    always @(spike_out_source_array[215]) begin 
        spike_out_source215 = spike_out_source_array[215];
    end
    always @(spike_out_source_array[216]) begin 
        spike_out_source216 = spike_out_source_array[216];
    end
    always @(spike_out_source_array[217]) begin 
        spike_out_source217 = spike_out_source_array[217];
    end
    always @(spike_out_source_array[218]) begin 
        spike_out_source218 = spike_out_source_array[218];
    end
    always @(spike_out_source_array[219]) begin 
        spike_out_source219 = spike_out_source_array[219];
    end
    always @(spike_out_source_array[220]) begin 
        spike_out_source220 = spike_out_source_array[220];
    end
    always @(spike_out_source_array[221]) begin 
        spike_out_source221 = spike_out_source_array[221];
    end
    always @(spike_out_source_array[222]) begin 
        spike_out_source222 = spike_out_source_array[222];
    end
    always @(spike_out_source_array[223]) begin 
        spike_out_source223 = spike_out_source_array[223];
    end
    always @(spike_out_source_array[224]) begin 
        spike_out_source224 = spike_out_source_array[224];
    end
    always @(spike_out_source_array[225]) begin 
        spike_out_source225 = spike_out_source_array[225];
    end
    always @(spike_out_source_array[226]) begin 
        spike_out_source226 = spike_out_source_array[226];
    end
    always @(spike_out_source_array[227]) begin 
        spike_out_source227 = spike_out_source_array[227];
    end
    always @(spike_out_source_array[228]) begin 
        spike_out_source228 = spike_out_source_array[228];
    end
    always @(spike_out_source_array[229]) begin 
        spike_out_source229 = spike_out_source_array[229];
    end
    always @(spike_out_source_array[230]) begin 
        spike_out_source230 = spike_out_source_array[230];
    end
    always @(spike_out_source_array[231]) begin 
        spike_out_source231 = spike_out_source_array[231];
    end
    always @(spike_out_source_array[232]) begin 
        spike_out_source232 = spike_out_source_array[232];
    end
    always @(spike_out_source_array[233]) begin 
        spike_out_source233 = spike_out_source_array[233];
    end
    always @(spike_out_source_array[234]) begin 
        spike_out_source234 = spike_out_source_array[234];
    end
    always @(spike_out_source_array[235]) begin 
        spike_out_source235 = spike_out_source_array[235];
    end
    always @(spike_out_source_array[236]) begin 
        spike_out_source236 = spike_out_source_array[236];
    end
    always @(spike_out_source_array[237]) begin 
        spike_out_source237 = spike_out_source_array[237];
    end
    always @(spike_out_source_array[238]) begin 
        spike_out_source238 = spike_out_source_array[238];
    end
    always @(spike_out_source_array[239]) begin 
        spike_out_source239 = spike_out_source_array[239];
    end
    always @(spike_out_source_array[240]) begin 
        spike_out_source240 = spike_out_source_array[240];
    end
    always @(spike_out_source_array[241]) begin 
        spike_out_source241 = spike_out_source_array[241];
    end
    always @(spike_out_source_array[242]) begin 
        spike_out_source242 = spike_out_source_array[242];
    end
    always @(spike_out_source_array[243]) begin 
        spike_out_source243 = spike_out_source_array[243];
    end
    always @(spike_out_source_array[244]) begin 
        spike_out_source244 = spike_out_source_array[244];
    end
    always @(spike_out_source_array[245]) begin 
        spike_out_source245 = spike_out_source_array[245];
    end
    always @(spike_out_source_array[246]) begin 
        spike_out_source246 = spike_out_source_array[246];
    end
    always @(spike_out_source_array[247]) begin 
        spike_out_source247 = spike_out_source_array[247];
    end
    always @(spike_out_source_array[248]) begin 
        spike_out_source248 = spike_out_source_array[248];
    end
    always @(spike_out_source_array[249]) begin 
        spike_out_source249 = spike_out_source_array[249];
    end
    always @(spike_out_source_array[250]) begin 
        spike_out_source250 = spike_out_source_array[250];
    end
    always @(spike_out_source_array[251]) begin 
        spike_out_source251 = spike_out_source_array[251];
    end
    always @(spike_out_source_array[252]) begin 
        spike_out_source252 = spike_out_source_array[252];
    end
    always @(spike_out_source_array[253]) begin 
        spike_out_source253 = spike_out_source_array[253];
    end
    always @(spike_out_source_array[254]) begin 
        spike_out_source254 = spike_out_source_array[254];
    end
    always @(spike_out_source_array[255]) begin 
        spike_out_source255 = spike_out_source_array[255];
    end
    always @(spike_out_source_array[256]) begin 
        spike_out_source256 = spike_out_source_array[256];
    end
    always @(spike_out_source_array[257]) begin 
        spike_out_source257 = spike_out_source_array[257];
    end
    always @(spike_out_source_array[258]) begin 
        spike_out_source258 = spike_out_source_array[258];
    end
    always @(spike_out_source_array[259]) begin 
        spike_out_source259 = spike_out_source_array[259];
    end
    always @(spike_out_source_array[260]) begin 
        spike_out_source260 = spike_out_source_array[260];
    end
    always @(spike_out_source_array[261]) begin 
        spike_out_source261 = spike_out_source_array[261];
    end
    always @(spike_out_source_array[262]) begin 
        spike_out_source262 = spike_out_source_array[262];
    end
    always @(spike_out_source_array[263]) begin 
        spike_out_source263 = spike_out_source_array[263];
    end
    always @(spike_out_source_array[264]) begin 
        spike_out_source264 = spike_out_source_array[264];
    end
    always @(spike_out_source_array[265]) begin 
        spike_out_source265 = spike_out_source_array[265];
    end
    always @(spike_out_source_array[266]) begin 
        spike_out_source266 = spike_out_source_array[266];
    end
    always @(spike_out_source_array[267]) begin 
        spike_out_source267 = spike_out_source_array[267];
    end
    always @(spike_out_source_array[268]) begin 
        spike_out_source268 = spike_out_source_array[268];
    end
    always @(spike_out_source_array[269]) begin 
        spike_out_source269 = spike_out_source_array[269];
    end
    always @(spike_out_source_array[270]) begin 
        spike_out_source270 = spike_out_source_array[270];
    end
    always @(spike_out_source_array[271]) begin 
        spike_out_source271 = spike_out_source_array[271];
    end
    always @(spike_out_source_array[272]) begin 
        spike_out_source272 = spike_out_source_array[272];
    end
    always @(spike_out_source_array[273]) begin 
        spike_out_source273 = spike_out_source_array[273];
    end
    always @(spike_out_source_array[274]) begin 
        spike_out_source274 = spike_out_source_array[274];
    end
    always @(spike_out_source_array[275]) begin 
        spike_out_source275 = spike_out_source_array[275];
    end
    always @(spike_out_source_array[276]) begin 
        spike_out_source276 = spike_out_source_array[276];
    end
    always @(spike_out_source_array[277]) begin 
        spike_out_source277 = spike_out_source_array[277];
    end
    always @(spike_out_source_array[278]) begin 
        spike_out_source278 = spike_out_source_array[278];
    end
    always @(spike_out_source_array[279]) begin 
        spike_out_source279 = spike_out_source_array[279];
    end
    always @(spike_out_source_array[280]) begin 
        spike_out_source280 = spike_out_source_array[280];
    end
    always @(spike_out_source_array[281]) begin 
        spike_out_source281 = spike_out_source_array[281];
    end
    always @(spike_out_source_array[282]) begin 
        spike_out_source282 = spike_out_source_array[282];
    end
    always @(spike_out_source_array[283]) begin 
        spike_out_source283 = spike_out_source_array[283];
    end
    always @(spike_out_source_array[284]) begin 
        spike_out_source284 = spike_out_source_array[284];
    end
    always @(spike_out_source_array[285]) begin 
        spike_out_source285 = spike_out_source_array[285];
    end
    always @(spike_out_source_array[286]) begin 
        spike_out_source286 = spike_out_source_array[286];
    end
    always @(spike_out_source_array[287]) begin 
        spike_out_source287 = spike_out_source_array[287];
    end
    always @(spike_out_source_array[288]) begin 
        spike_out_source288 = spike_out_source_array[288];
    end
    always @(spike_out_source_array[289]) begin 
        spike_out_source289 = spike_out_source_array[289];
    end
    always @(spike_out_source_array[290]) begin 
        spike_out_source290 = spike_out_source_array[290];
    end
    always @(spike_out_source_array[291]) begin 
        spike_out_source291 = spike_out_source_array[291];
    end
    always @(spike_out_source_array[292]) begin 
        spike_out_source292 = spike_out_source_array[292];
    end
    always @(spike_out_source_array[293]) begin 
        spike_out_source293 = spike_out_source_array[293];
    end
    always @(spike_out_source_array[294]) begin 
        spike_out_source294 = spike_out_source_array[294];
    end
    always @(spike_out_source_array[295]) begin 
        spike_out_source295 = spike_out_source_array[295];
    end
    always @(spike_out_source_array[296]) begin 
        spike_out_source296 = spike_out_source_array[296];
    end
    always @(spike_out_source_array[297]) begin 
        spike_out_source297 = spike_out_source_array[297];
    end
    always @(spike_out_source_array[298]) begin 
        spike_out_source298 = spike_out_source_array[298];
    end
    always @(spike_out_source_array[299]) begin 
        spike_out_source299 = spike_out_source_array[299];
    end
    always @(spike_out_source_array[300]) begin 
        spike_out_source300 = spike_out_source_array[300];
    end
    always @(spike_out_source_array[301]) begin 
        spike_out_source301 = spike_out_source_array[301];
    end
    always @(spike_out_source_array[302]) begin 
        spike_out_source302 = spike_out_source_array[302];
    end
    always @(spike_out_source_array[303]) begin 
        spike_out_source303 = spike_out_source_array[303];
    end
    always @(spike_out_source_array[304]) begin 
        spike_out_source304 = spike_out_source_array[304];
    end
    always @(spike_out_source_array[305]) begin 
        spike_out_source305 = spike_out_source_array[305];
    end
    always @(spike_out_source_array[306]) begin 
        spike_out_source306 = spike_out_source_array[306];
    end
    always @(spike_out_source_array[307]) begin 
        spike_out_source307 = spike_out_source_array[307];
    end
    always @(spike_out_source_array[308]) begin 
        spike_out_source308 = spike_out_source_array[308];
    end
    always @(spike_out_source_array[309]) begin 
        spike_out_source309 = spike_out_source_array[309];
    end
    always @(spike_out_source_array[310]) begin 
        spike_out_source310 = spike_out_source_array[310];
    end
    always @(spike_out_source_array[311]) begin 
        spike_out_source311 = spike_out_source_array[311];
    end
    always @(spike_out_source_array[312]) begin 
        spike_out_source312 = spike_out_source_array[312];
    end
    always @(spike_out_source_array[313]) begin 
        spike_out_source313 = spike_out_source_array[313];
    end
    always @(spike_out_source_array[314]) begin 
        spike_out_source314 = spike_out_source_array[314];
    end
    always @(spike_out_source_array[315]) begin 
        spike_out_source315 = spike_out_source_array[315];
    end
    always @(spike_out_source_array[316]) begin 
        spike_out_source316 = spike_out_source_array[316];
    end
    always @(spike_out_source_array[317]) begin 
        spike_out_source317 = spike_out_source_array[317];
    end
    always @(spike_out_source_array[318]) begin 
        spike_out_source318 = spike_out_source_array[318];
    end
    always @(spike_out_source_array[319]) begin 
        spike_out_source319 = spike_out_source_array[319];
    end
    always @(spike_out_source_array[320]) begin 
        spike_out_source320 = spike_out_source_array[320];
    end
    always @(spike_out_source_array[321]) begin 
        spike_out_source321 = spike_out_source_array[321];
    end
    always @(spike_out_source_array[322]) begin 
        spike_out_source322 = spike_out_source_array[322];
    end
    always @(spike_out_source_array[323]) begin 
        spike_out_source323 = spike_out_source_array[323];
    end
    always @(spike_out_source_array[324]) begin 
        spike_out_source324 = spike_out_source_array[324];
    end
    always @(spike_out_source_array[325]) begin 
        spike_out_source325 = spike_out_source_array[325];
    end
    always @(spike_out_source_array[326]) begin 
        spike_out_source326 = spike_out_source_array[326];
    end
    always @(spike_out_source_array[327]) begin 
        spike_out_source327 = spike_out_source_array[327];
    end
    always @(spike_out_source_array[328]) begin 
        spike_out_source328 = spike_out_source_array[328];
    end
    always @(spike_out_source_array[329]) begin 
        spike_out_source329 = spike_out_source_array[329];
    end
    always @(spike_out_source_array[330]) begin 
        spike_out_source330 = spike_out_source_array[330];
    end
    always @(spike_out_source_array[331]) begin 
        spike_out_source331 = spike_out_source_array[331];
    end
    always @(spike_out_source_array[332]) begin 
        spike_out_source332 = spike_out_source_array[332];
    end
    always @(spike_out_source_array[333]) begin 
        spike_out_source333 = spike_out_source_array[333];
    end
    always @(spike_out_source_array[334]) begin 
        spike_out_source334 = spike_out_source_array[334];
    end
    always @(spike_out_source_array[335]) begin 
        spike_out_source335 = spike_out_source_array[335];
    end
    always @(spike_out_source_array[336]) begin 
        spike_out_source336 = spike_out_source_array[336];
    end
    always @(spike_out_source_array[337]) begin 
        spike_out_source337 = spike_out_source_array[337];
    end
    always @(spike_out_source_array[338]) begin 
        spike_out_source338 = spike_out_source_array[338];
    end
    always @(spike_out_source_array[339]) begin 
        spike_out_source339 = spike_out_source_array[339];
    end
    always @(spike_out_source_array[340]) begin 
        spike_out_source340 = spike_out_source_array[340];
    end
    always @(spike_out_source_array[341]) begin 
        spike_out_source341 = spike_out_source_array[341];
    end
    always @(spike_out_source_array[342]) begin 
        spike_out_source342 = spike_out_source_array[342];
    end
    always @(spike_out_source_array[343]) begin 
        spike_out_source343 = spike_out_source_array[343];
    end
    always @(spike_out_source_array[344]) begin 
        spike_out_source344 = spike_out_source_array[344];
    end
    always @(spike_out_source_array[345]) begin 
        spike_out_source345 = spike_out_source_array[345];
    end
    always @(spike_out_source_array[346]) begin 
        spike_out_source346 = spike_out_source_array[346];
    end
    always @(spike_out_source_array[347]) begin 
        spike_out_source347 = spike_out_source_array[347];
    end
    always @(spike_out_source_array[348]) begin 
        spike_out_source348 = spike_out_source_array[348];
    end
    always @(spike_out_source_array[349]) begin 
        spike_out_source349 = spike_out_source_array[349];
    end
    always @(spike_out_source_array[350]) begin 
        spike_out_source350 = spike_out_source_array[350];
    end
    always @(spike_out_source_array[351]) begin 
        spike_out_source351 = spike_out_source_array[351];
    end
    always @(spike_out_source_array[352]) begin 
        spike_out_source352 = spike_out_source_array[352];
    end
    always @(spike_out_source_array[353]) begin 
        spike_out_source353 = spike_out_source_array[353];
    end
    always @(spike_out_source_array[354]) begin 
        spike_out_source354 = spike_out_source_array[354];
    end
    always @(spike_out_source_array[355]) begin 
        spike_out_source355 = spike_out_source_array[355];
    end
    always @(spike_out_source_array[356]) begin 
        spike_out_source356 = spike_out_source_array[356];
    end
    always @(spike_out_source_array[357]) begin 
        spike_out_source357 = spike_out_source_array[357];
    end
    always @(spike_out_source_array[358]) begin 
        spike_out_source358 = spike_out_source_array[358];
    end
    always @(spike_out_source_array[359]) begin 
        spike_out_source359 = spike_out_source_array[359];
    end
    always @(spike_out_source_array[360]) begin 
        spike_out_source360 = spike_out_source_array[360];
    end
    always @(spike_out_source_array[361]) begin 
        spike_out_source361 = spike_out_source_array[361];
    end
    always @(spike_out_source_array[362]) begin 
        spike_out_source362 = spike_out_source_array[362];
    end
    always @(spike_out_source_array[363]) begin 
        spike_out_source363 = spike_out_source_array[363];
    end
    always @(spike_out_source_array[364]) begin 
        spike_out_source364 = spike_out_source_array[364];
    end
    always @(spike_out_source_array[365]) begin 
        spike_out_source365 = spike_out_source_array[365];
    end
    always @(spike_out_source_array[366]) begin 
        spike_out_source366 = spike_out_source_array[366];
    end
    always @(spike_out_source_array[367]) begin 
        spike_out_source367 = spike_out_source_array[367];
    end
    always @(spike_out_source_array[368]) begin 
        spike_out_source368 = spike_out_source_array[368];
    end
    always @(spike_out_source_array[369]) begin 
        spike_out_source369 = spike_out_source_array[369];
    end
    always @(spike_out_source_array[370]) begin 
        spike_out_source370 = spike_out_source_array[370];
    end
    always @(spike_out_source_array[371]) begin 
        spike_out_source371 = spike_out_source_array[371];
    end
    always @(spike_out_source_array[372]) begin 
        spike_out_source372 = spike_out_source_array[372];
    end
    always @(spike_out_source_array[373]) begin 
        spike_out_source373 = spike_out_source_array[373];
    end
    always @(spike_out_source_array[374]) begin 
        spike_out_source374 = spike_out_source_array[374];
    end
    always @(spike_out_source_array[375]) begin 
        spike_out_source375 = spike_out_source_array[375];
    end
    always @(spike_out_source_array[376]) begin 
        spike_out_source376 = spike_out_source_array[376];
    end
    always @(spike_out_source_array[377]) begin 
        spike_out_source377 = spike_out_source_array[377];
    end
    always @(spike_out_source_array[378]) begin 
        spike_out_source378 = spike_out_source_array[378];
    end
    always @(spike_out_source_array[379]) begin 
        spike_out_source379 = spike_out_source_array[379];
    end
    always @(spike_out_source_array[380]) begin 
        spike_out_source380 = spike_out_source_array[380];
    end
    always @(spike_out_source_array[381]) begin 
        spike_out_source381 = spike_out_source_array[381];
    end
    always @(spike_out_source_array[382]) begin 
        spike_out_source382 = spike_out_source_array[382];
    end
    always @(spike_out_source_array[383]) begin 
        spike_out_source383 = spike_out_source_array[383];
    end
    always @(spike_out_source_array[384]) begin 
        spike_out_source384 = spike_out_source_array[384];
    end
    always @(spike_out_source_array[385]) begin 
        spike_out_source385 = spike_out_source_array[385];
    end
    always @(spike_out_source_array[386]) begin 
        spike_out_source386 = spike_out_source_array[386];
    end
    always @(spike_out_source_array[387]) begin 
        spike_out_source387 = spike_out_source_array[387];
    end
    always @(spike_out_source_array[388]) begin 
        spike_out_source388 = spike_out_source_array[388];
    end
    always @(spike_out_source_array[389]) begin 
        spike_out_source389 = spike_out_source_array[389];
    end
    always @(spike_out_source_array[390]) begin 
        spike_out_source390 = spike_out_source_array[390];
    end
    always @(spike_out_source_array[391]) begin 
        spike_out_source391 = spike_out_source_array[391];
    end
    always @(spike_out_source_array[392]) begin 
        spike_out_source392 = spike_out_source_array[392];
    end
    always @(spike_out_source_array[393]) begin 
        spike_out_source393 = spike_out_source_array[393];
    end
    always @(spike_out_source_array[394]) begin 
        spike_out_source394 = spike_out_source_array[394];
    end
    always @(spike_out_source_array[395]) begin 
        spike_out_source395 = spike_out_source_array[395];
    end
    always @(spike_out_source_array[396]) begin 
        spike_out_source396 = spike_out_source_array[396];
    end
    always @(spike_out_source_array[397]) begin 
        spike_out_source397 = spike_out_source_array[397];
    end
    always @(spike_out_source_array[398]) begin 
        spike_out_source398 = spike_out_source_array[398];
    end
    always @(spike_out_source_array[399]) begin 
        spike_out_source399 = spike_out_source_array[399];
    end
    always @(spike_out_source_array[400]) begin 
        spike_out_source400 = spike_out_source_array[400];
    end
    always @(spike_out_source_array[401]) begin 
        spike_out_source401 = spike_out_source_array[401];
    end
    always @(spike_out_source_array[402]) begin 
        spike_out_source402 = spike_out_source_array[402];
    end
    always @(spike_out_source_array[403]) begin 
        spike_out_source403 = spike_out_source_array[403];
    end
    always @(spike_out_source_array[404]) begin 
        spike_out_source404 = spike_out_source_array[404];
    end
    always @(spike_out_source_array[405]) begin 
        spike_out_source405 = spike_out_source_array[405];
    end
    always @(spike_out_source_array[406]) begin 
        spike_out_source406 = spike_out_source_array[406];
    end
    always @(spike_out_source_array[407]) begin 
        spike_out_source407 = spike_out_source_array[407];
    end
    always @(spike_out_source_array[408]) begin 
        spike_out_source408 = spike_out_source_array[408];
    end
    always @(spike_out_source_array[409]) begin 
        spike_out_source409 = spike_out_source_array[409];
    end
    always @(spike_out_source_array[410]) begin 
        spike_out_source410 = spike_out_source_array[410];
    end
    always @(spike_out_source_array[411]) begin 
        spike_out_source411 = spike_out_source_array[411];
    end
    always @(spike_out_source_array[412]) begin 
        spike_out_source412 = spike_out_source_array[412];
    end
    always @(spike_out_source_array[413]) begin 
        spike_out_source413 = spike_out_source_array[413];
    end
    always @(spike_out_source_array[414]) begin 
        spike_out_source414 = spike_out_source_array[414];
    end
    always @(spike_out_source_array[415]) begin 
        spike_out_source415 = spike_out_source_array[415];
    end
    always @(spike_out_source_array[416]) begin 
        spike_out_source416 = spike_out_source_array[416];
    end
    always @(spike_out_source_array[417]) begin 
        spike_out_source417 = spike_out_source_array[417];
    end
    always @(spike_out_source_array[418]) begin 
        spike_out_source418 = spike_out_source_array[418];
    end
    always @(spike_out_source_array[419]) begin 
        spike_out_source419 = spike_out_source_array[419];
    end
    always @(spike_out_source_array[420]) begin 
        spike_out_source420 = spike_out_source_array[420];
    end
    always @(spike_out_source_array[421]) begin 
        spike_out_source421 = spike_out_source_array[421];
    end
    always @(spike_out_source_array[422]) begin 
        spike_out_source422 = spike_out_source_array[422];
    end
    always @(spike_out_source_array[423]) begin 
        spike_out_source423 = spike_out_source_array[423];
    end
    always @(spike_out_source_array[424]) begin 
        spike_out_source424 = spike_out_source_array[424];
    end
    always @(spike_out_source_array[425]) begin 
        spike_out_source425 = spike_out_source_array[425];
    end
    always @(spike_out_source_array[426]) begin 
        spike_out_source426 = spike_out_source_array[426];
    end
    always @(spike_out_source_array[427]) begin 
        spike_out_source427 = spike_out_source_array[427];
    end
    always @(spike_out_source_array[428]) begin 
        spike_out_source428 = spike_out_source_array[428];
    end
    always @(spike_out_source_array[429]) begin 
        spike_out_source429 = spike_out_source_array[429];
    end
    always @(spike_out_source_array[430]) begin 
        spike_out_source430 = spike_out_source_array[430];
    end
    always @(spike_out_source_array[431]) begin 
        spike_out_source431 = spike_out_source_array[431];
    end
    always @(spike_out_source_array[432]) begin 
        spike_out_source432 = spike_out_source_array[432];
    end
    always @(spike_out_source_array[433]) begin 
        spike_out_source433 = spike_out_source_array[433];
    end
    always @(spike_out_source_array[434]) begin 
        spike_out_source434 = spike_out_source_array[434];
    end
    always @(spike_out_source_array[435]) begin 
        spike_out_source435 = spike_out_source_array[435];
    end
    always @(spike_out_source_array[436]) begin 
        spike_out_source436 = spike_out_source_array[436];
    end
    always @(spike_out_source_array[437]) begin 
        spike_out_source437 = spike_out_source_array[437];
    end
    always @(spike_out_source_array[438]) begin 
        spike_out_source438 = spike_out_source_array[438];
    end
    always @(spike_out_source_array[439]) begin 
        spike_out_source439 = spike_out_source_array[439];
    end
    always @(spike_out_source_array[440]) begin 
        spike_out_source440 = spike_out_source_array[440];
    end
    always @(spike_out_source_array[441]) begin 
        spike_out_source441 = spike_out_source_array[441];
    end
    always @(spike_out_source_array[442]) begin 
        spike_out_source442 = spike_out_source_array[442];
    end
    always @(spike_out_source_array[443]) begin 
        spike_out_source443 = spike_out_source_array[443];
    end
    always @(spike_out_source_array[444]) begin 
        spike_out_source444 = spike_out_source_array[444];
    end
    always @(spike_out_source_array[445]) begin 
        spike_out_source445 = spike_out_source_array[445];
    end
    always @(spike_out_source_array[446]) begin 
        spike_out_source446 = spike_out_source_array[446];
    end
    always @(spike_out_source_array[447]) begin 
        spike_out_source447 = spike_out_source_array[447];
    end
    always @(spike_out_source_array[448]) begin 
        spike_out_source448 = spike_out_source_array[448];
    end
    always @(spike_out_source_array[449]) begin 
        spike_out_source449 = spike_out_source_array[449];
    end
    always @(spike_out_source_array[450]) begin 
        spike_out_source450 = spike_out_source_array[450];
    end
    always @(spike_out_source_array[451]) begin 
        spike_out_source451 = spike_out_source_array[451];
    end
    always @(spike_out_source_array[452]) begin 
        spike_out_source452 = spike_out_source_array[452];
    end
    always @(spike_out_source_array[453]) begin 
        spike_out_source453 = spike_out_source_array[453];
    end
    always @(spike_out_source_array[454]) begin 
        spike_out_source454 = spike_out_source_array[454];
    end
    always @(spike_out_source_array[455]) begin 
        spike_out_source455 = spike_out_source_array[455];
    end
    always @(spike_out_source_array[456]) begin 
        spike_out_source456 = spike_out_source_array[456];
    end
    always @(spike_out_source_array[457]) begin 
        spike_out_source457 = spike_out_source_array[457];
    end
    always @(spike_out_source_array[458]) begin 
        spike_out_source458 = spike_out_source_array[458];
    end
    always @(spike_out_source_array[459]) begin 
        spike_out_source459 = spike_out_source_array[459];
    end
    always @(spike_out_source_array[460]) begin 
        spike_out_source460 = spike_out_source_array[460];
    end
    always @(spike_out_source_array[461]) begin 
        spike_out_source461 = spike_out_source_array[461];
    end
    always @(spike_out_source_array[462]) begin 
        spike_out_source462 = spike_out_source_array[462];
    end
    always @(spike_out_source_array[463]) begin 
        spike_out_source463 = spike_out_source_array[463];
    end
    always @(spike_out_source_array[464]) begin 
        spike_out_source464 = spike_out_source_array[464];
    end
    always @(spike_out_source_array[465]) begin 
        spike_out_source465 = spike_out_source_array[465];
    end
    always @(spike_out_source_array[466]) begin 
        spike_out_source466 = spike_out_source_array[466];
    end
    always @(spike_out_source_array[467]) begin 
        spike_out_source467 = spike_out_source_array[467];
    end
    always @(spike_out_source_array[468]) begin 
        spike_out_source468 = spike_out_source_array[468];
    end
    always @(spike_out_source_array[469]) begin 
        spike_out_source469 = spike_out_source_array[469];
    end
    always @(spike_out_source_array[470]) begin 
        spike_out_source470 = spike_out_source_array[470];
    end
    always @(spike_out_source_array[471]) begin 
        spike_out_source471 = spike_out_source_array[471];
    end
    always @(spike_out_source_array[472]) begin 
        spike_out_source472 = spike_out_source_array[472];
    end
    always @(spike_out_source_array[473]) begin 
        spike_out_source473 = spike_out_source_array[473];
    end
    always @(spike_out_source_array[474]) begin 
        spike_out_source474 = spike_out_source_array[474];
    end
    always @(spike_out_source_array[475]) begin 
        spike_out_source475 = spike_out_source_array[475];
    end
    always @(spike_out_source_array[476]) begin 
        spike_out_source476 = spike_out_source_array[476];
    end
    always @(spike_out_source_array[477]) begin 
        spike_out_source477 = spike_out_source_array[477];
    end
    always @(spike_out_source_array[478]) begin 
        spike_out_source478 = spike_out_source_array[478];
    end
    always @(spike_out_source_array[479]) begin 
        spike_out_source479 = spike_out_source_array[479];
    end
    always @(spike_out_source_array[480]) begin 
        spike_out_source480 = spike_out_source_array[480];
    end
    always @(spike_out_source_array[481]) begin 
        spike_out_source481 = spike_out_source_array[481];
    end
    always @(spike_out_source_array[482]) begin 
        spike_out_source482 = spike_out_source_array[482];
    end
    always @(spike_out_source_array[483]) begin 
        spike_out_source483 = spike_out_source_array[483];
    end
    always @(spike_out_source_array[484]) begin 
        spike_out_source484 = spike_out_source_array[484];
    end
    always @(spike_out_source_array[485]) begin 
        spike_out_source485 = spike_out_source_array[485];
    end
    always @(spike_out_source_array[486]) begin 
        spike_out_source486 = spike_out_source_array[486];
    end
    always @(spike_out_source_array[487]) begin 
        spike_out_source487 = spike_out_source_array[487];
    end
    always @(spike_out_source_array[488]) begin 
        spike_out_source488 = spike_out_source_array[488];
    end
    always @(spike_out_source_array[489]) begin 
        spike_out_source489 = spike_out_source_array[489];
    end
    always @(spike_out_source_array[490]) begin 
        spike_out_source490 = spike_out_source_array[490];
    end
    always @(spike_out_source_array[491]) begin 
        spike_out_source491 = spike_out_source_array[491];
    end
    always @(spike_out_source_array[492]) begin 
        spike_out_source492 = spike_out_source_array[492];
    end
    always @(spike_out_source_array[493]) begin 
        spike_out_source493 = spike_out_source_array[493];
    end
    always @(spike_out_source_array[494]) begin 
        spike_out_source494 = spike_out_source_array[494];
    end
    always @(spike_out_source_array[495]) begin 
        spike_out_source495 = spike_out_source_array[495];
    end
    always @(spike_out_source_array[496]) begin 
        spike_out_source496 = spike_out_source_array[496];
    end
    always @(spike_out_source_array[497]) begin 
        spike_out_source497 = spike_out_source_array[497];
    end
    always @(spike_out_source_array[498]) begin 
        spike_out_source498 = spike_out_source_array[498];
    end
    always @(spike_out_source_array[499]) begin 
        spike_out_source499 = spike_out_source_array[499];
    end
    always @(spike_out_source_array[500]) begin 
        spike_out_source500 = spike_out_source_array[500];
    end
    always @(spike_out_source_array[501]) begin 
        spike_out_source501 = spike_out_source_array[501];
    end
    always @(spike_out_source_array[502]) begin 
        spike_out_source502 = spike_out_source_array[502];
    end
    always @(spike_out_source_array[503]) begin 
        spike_out_source503 = spike_out_source_array[503];
    end
    always @(spike_out_source_array[504]) begin 
        spike_out_source504 = spike_out_source_array[504];
    end
    always @(spike_out_source_array[505]) begin 
        spike_out_source505 = spike_out_source_array[505];
    end
    always @(spike_out_source_array[506]) begin 
        spike_out_source506 = spike_out_source_array[506];
    end
    always @(spike_out_source_array[507]) begin 
        spike_out_source507 = spike_out_source_array[507];
    end
    always @(spike_out_source_array[508]) begin 
        spike_out_source508 = spike_out_source_array[508];
    end
    always @(spike_out_source_array[509]) begin 
        spike_out_source509 = spike_out_source_array[509];
    end
    always @(spike_out_source_array[510]) begin 
        spike_out_source510 = spike_out_source_array[510];
    end
    always @(spike_out_source_array[511]) begin 
        spike_out_source511 = spike_out_source_array[511];
    end
    always @(spike_out_source_array[512]) begin 
        spike_out_source512 = spike_out_source_array[512];
    end
    always @(spike_out_source_array[513]) begin 
        spike_out_source513 = spike_out_source_array[513];
    end
    always @(spike_out_source_array[514]) begin 
        spike_out_source514 = spike_out_source_array[514];
    end
    always @(spike_out_source_array[515]) begin 
        spike_out_source515 = spike_out_source_array[515];
    end
    always @(spike_out_source_array[516]) begin 
        spike_out_source516 = spike_out_source_array[516];
    end
    always @(spike_out_source_array[517]) begin 
        spike_out_source517 = spike_out_source_array[517];
    end
    always @(spike_out_source_array[518]) begin 
        spike_out_source518 = spike_out_source_array[518];
    end
    always @(spike_out_source_array[519]) begin 
        spike_out_source519 = spike_out_source_array[519];
    end
    always @(spike_out_source_array[520]) begin 
        spike_out_source520 = spike_out_source_array[520];
    end
    always @(spike_out_source_array[521]) begin 
        spike_out_source521 = spike_out_source_array[521];
    end
    always @(spike_out_source_array[522]) begin 
        spike_out_source522 = spike_out_source_array[522];
    end
    always @(spike_out_source_array[523]) begin 
        spike_out_source523 = spike_out_source_array[523];
    end
    always @(spike_out_source_array[524]) begin 
        spike_out_source524 = spike_out_source_array[524];
    end
    always @(spike_out_source_array[525]) begin 
        spike_out_source525 = spike_out_source_array[525];
    end
    always @(spike_out_source_array[526]) begin 
        spike_out_source526 = spike_out_source_array[526];
    end
    always @(spike_out_source_array[527]) begin 
        spike_out_source527 = spike_out_source_array[527];
    end
    always @(spike_out_source_array[528]) begin 
        spike_out_source528 = spike_out_source_array[528];
    end
    always @(spike_out_source_array[529]) begin 
        spike_out_source529 = spike_out_source_array[529];
    end
    always @(spike_out_source_array[530]) begin 
        spike_out_source530 = spike_out_source_array[530];
    end
    always @(spike_out_source_array[531]) begin 
        spike_out_source531 = spike_out_source_array[531];
    end
    always @(spike_out_source_array[532]) begin 
        spike_out_source532 = spike_out_source_array[532];
    end
    always @(spike_out_source_array[533]) begin 
        spike_out_source533 = spike_out_source_array[533];
    end
    always @(spike_out_source_array[534]) begin 
        spike_out_source534 = spike_out_source_array[534];
    end
    always @(spike_out_source_array[535]) begin 
        spike_out_source535 = spike_out_source_array[535];
    end
    always @(spike_out_source_array[536]) begin 
        spike_out_source536 = spike_out_source_array[536];
    end
    always @(spike_out_source_array[537]) begin 
        spike_out_source537 = spike_out_source_array[537];
    end
    always @(spike_out_source_array[538]) begin 
        spike_out_source538 = spike_out_source_array[538];
    end
    always @(spike_out_source_array[539]) begin 
        spike_out_source539 = spike_out_source_array[539];
    end
    always @(spike_out_source_array[540]) begin 
        spike_out_source540 = spike_out_source_array[540];
    end
    always @(spike_out_source_array[541]) begin 
        spike_out_source541 = spike_out_source_array[541];
    end
    always @(spike_out_source_array[542]) begin 
        spike_out_source542 = spike_out_source_array[542];
    end
    always @(spike_out_source_array[543]) begin 
        spike_out_source543 = spike_out_source_array[543];
    end
    always @(spike_out_source_array[544]) begin 
        spike_out_source544 = spike_out_source_array[544];
    end
    always @(spike_out_source_array[545]) begin 
        spike_out_source545 = spike_out_source_array[545];
    end
    always @(spike_out_source_array[546]) begin 
        spike_out_source546 = spike_out_source_array[546];
    end
    always @(spike_out_source_array[547]) begin 
        spike_out_source547 = spike_out_source_array[547];
    end
    always @(spike_out_source_array[548]) begin 
        spike_out_source548 = spike_out_source_array[548];
    end
    always @(spike_out_source_array[549]) begin 
        spike_out_source549 = spike_out_source_array[549];
    end
    always @(spike_out_source_array[550]) begin 
        spike_out_source550 = spike_out_source_array[550];
    end
    always @(spike_out_source_array[551]) begin 
        spike_out_source551 = spike_out_source_array[551];
    end
    always @(spike_out_source_array[552]) begin 
        spike_out_source552 = spike_out_source_array[552];
    end
    always @(spike_out_source_array[553]) begin 
        spike_out_source553 = spike_out_source_array[553];
    end
    always @(spike_out_source_array[554]) begin 
        spike_out_source554 = spike_out_source_array[554];
    end
    always @(spike_out_source_array[555]) begin 
        spike_out_source555 = spike_out_source_array[555];
    end
    always @(spike_out_source_array[556]) begin 
        spike_out_source556 = spike_out_source_array[556];
    end
    always @(spike_out_source_array[557]) begin 
        spike_out_source557 = spike_out_source_array[557];
    end
    always @(spike_out_source_array[558]) begin 
        spike_out_source558 = spike_out_source_array[558];
    end
    always @(spike_out_source_array[559]) begin 
        spike_out_source559 = spike_out_source_array[559];
    end
    always @(spike_out_source_array[560]) begin 
        spike_out_source560 = spike_out_source_array[560];
    end
    always @(spike_out_source_array[561]) begin 
        spike_out_source561 = spike_out_source_array[561];
    end
    always @(spike_out_source_array[562]) begin 
        spike_out_source562 = spike_out_source_array[562];
    end
    always @(spike_out_source_array[563]) begin 
        spike_out_source563 = spike_out_source_array[563];
    end
    always @(spike_out_source_array[564]) begin 
        spike_out_source564 = spike_out_source_array[564];
    end
    always @(spike_out_source_array[565]) begin 
        spike_out_source565 = spike_out_source_array[565];
    end
    always @(spike_out_source_array[566]) begin 
        spike_out_source566 = spike_out_source_array[566];
    end
    always @(spike_out_source_array[567]) begin 
        spike_out_source567 = spike_out_source_array[567];
    end
    always @(spike_out_source_array[568]) begin 
        spike_out_source568 = spike_out_source_array[568];
    end
    always @(spike_out_source_array[569]) begin 
        spike_out_source569 = spike_out_source_array[569];
    end
    always @(spike_out_source_array[570]) begin 
        spike_out_source570 = spike_out_source_array[570];
    end
    always @(spike_out_source_array[571]) begin 
        spike_out_source571 = spike_out_source_array[571];
    end
    always @(spike_out_source_array[572]) begin 
        spike_out_source572 = spike_out_source_array[572];
    end
    always @(spike_out_source_array[573]) begin 
        spike_out_source573 = spike_out_source_array[573];
    end
    always @(spike_out_source_array[574]) begin 
        spike_out_source574 = spike_out_source_array[574];
    end
    always @(spike_out_source_array[575]) begin 
        spike_out_source575 = spike_out_source_array[575];
    end
    always @(spike_out_source_array[576]) begin 
        spike_out_source576 = spike_out_source_array[576];
    end
    always @(spike_out_source_array[577]) begin 
        spike_out_source577 = spike_out_source_array[577];
    end
    always @(spike_out_source_array[578]) begin 
        spike_out_source578 = spike_out_source_array[578];
    end
    always @(spike_out_source_array[579]) begin 
        spike_out_source579 = spike_out_source_array[579];
    end
    always @(spike_out_source_array[580]) begin 
        spike_out_source580 = spike_out_source_array[580];
    end
    always @(spike_out_source_array[581]) begin 
        spike_out_source581 = spike_out_source_array[581];
    end
    always @(spike_out_source_array[582]) begin 
        spike_out_source582 = spike_out_source_array[582];
    end
    always @(spike_out_source_array[583]) begin 
        spike_out_source583 = spike_out_source_array[583];
    end
    always @(spike_out_source_array[584]) begin 
        spike_out_source584 = spike_out_source_array[584];
    end
    always @(spike_out_source_array[585]) begin 
        spike_out_source585 = spike_out_source_array[585];
    end
    always @(spike_out_source_array[586]) begin 
        spike_out_source586 = spike_out_source_array[586];
    end
    always @(spike_out_source_array[587]) begin 
        spike_out_source587 = spike_out_source_array[587];
    end
    always @(spike_out_source_array[588]) begin 
        spike_out_source588 = spike_out_source_array[588];
    end
    always @(spike_out_source_array[589]) begin 
        spike_out_source589 = spike_out_source_array[589];
    end
    always @(spike_out_source_array[590]) begin 
        spike_out_source590 = spike_out_source_array[590];
    end
    always @(spike_out_source_array[591]) begin 
        spike_out_source591 = spike_out_source_array[591];
    end
    always @(spike_out_source_array[592]) begin 
        spike_out_source592 = spike_out_source_array[592];
    end
    always @(spike_out_source_array[593]) begin 
        spike_out_source593 = spike_out_source_array[593];
    end
    always @(spike_out_source_array[594]) begin 
        spike_out_source594 = spike_out_source_array[594];
    end
    always @(spike_out_source_array[595]) begin 
        spike_out_source595 = spike_out_source_array[595];
    end
    always @(spike_out_source_array[596]) begin 
        spike_out_source596 = spike_out_source_array[596];
    end
    always @(spike_out_source_array[597]) begin 
        spike_out_source597 = spike_out_source_array[597];
    end
    always @(spike_out_source_array[598]) begin 
        spike_out_source598 = spike_out_source_array[598];
    end
    always @(spike_out_source_array[599]) begin 
        spike_out_source599 = spike_out_source_array[599];
    end
    always @(spike_out_source_array[600]) begin 
        spike_out_source600 = spike_out_source_array[600];
    end
    always @(spike_out_source_array[601]) begin 
        spike_out_source601 = spike_out_source_array[601];
    end
    always @(spike_out_source_array[602]) begin 
        spike_out_source602 = spike_out_source_array[602];
    end
    always @(spike_out_source_array[603]) begin 
        spike_out_source603 = spike_out_source_array[603];
    end
    always @(spike_out_source_array[604]) begin 
        spike_out_source604 = spike_out_source_array[604];
    end
    always @(spike_out_source_array[605]) begin 
        spike_out_source605 = spike_out_source_array[605];
    end
    always @(spike_out_source_array[606]) begin 
        spike_out_source606 = spike_out_source_array[606];
    end
    always @(spike_out_source_array[607]) begin 
        spike_out_source607 = spike_out_source_array[607];
    end
    always @(spike_out_source_array[608]) begin 
        spike_out_source608 = spike_out_source_array[608];
    end
    always @(spike_out_source_array[609]) begin 
        spike_out_source609 = spike_out_source_array[609];
    end
    always @(spike_out_source_array[610]) begin 
        spike_out_source610 = spike_out_source_array[610];
    end
    always @(spike_out_source_array[611]) begin 
        spike_out_source611 = spike_out_source_array[611];
    end
    always @(spike_out_source_array[612]) begin 
        spike_out_source612 = spike_out_source_array[612];
    end
    always @(spike_out_source_array[613]) begin 
        spike_out_source613 = spike_out_source_array[613];
    end
    always @(spike_out_source_array[614]) begin 
        spike_out_source614 = spike_out_source_array[614];
    end
    always @(spike_out_source_array[615]) begin 
        spike_out_source615 = spike_out_source_array[615];
    end
    always @(spike_out_source_array[616]) begin 
        spike_out_source616 = spike_out_source_array[616];
    end
    always @(spike_out_source_array[617]) begin 
        spike_out_source617 = spike_out_source_array[617];
    end
    always @(spike_out_source_array[618]) begin 
        spike_out_source618 = spike_out_source_array[618];
    end
    always @(spike_out_source_array[619]) begin 
        spike_out_source619 = spike_out_source_array[619];
    end
    always @(spike_out_source_array[620]) begin 
        spike_out_source620 = spike_out_source_array[620];
    end
    always @(spike_out_source_array[621]) begin 
        spike_out_source621 = spike_out_source_array[621];
    end
    always @(spike_out_source_array[622]) begin 
        spike_out_source622 = spike_out_source_array[622];
    end
    always @(spike_out_source_array[623]) begin 
        spike_out_source623 = spike_out_source_array[623];
    end
    always @(spike_out_source_array[624]) begin 
        spike_out_source624 = spike_out_source_array[624];
    end
    always @(spike_out_source_array[625]) begin 
        spike_out_source625 = spike_out_source_array[625];
    end
    always @(spike_out_source_array[626]) begin 
        spike_out_source626 = spike_out_source_array[626];
    end
    always @(spike_out_source_array[627]) begin 
        spike_out_source627 = spike_out_source_array[627];
    end
    always @(spike_out_source_array[628]) begin 
        spike_out_source628 = spike_out_source_array[628];
    end
    always @(spike_out_source_array[629]) begin 
        spike_out_source629 = spike_out_source_array[629];
    end
    always @(spike_out_source_array[630]) begin 
        spike_out_source630 = spike_out_source_array[630];
    end
    always @(spike_out_source_array[631]) begin 
        spike_out_source631 = spike_out_source_array[631];
    end
    always @(spike_out_source_array[632]) begin 
        spike_out_source632 = spike_out_source_array[632];
    end
    always @(spike_out_source_array[633]) begin 
        spike_out_source633 = spike_out_source_array[633];
    end
    always @(spike_out_source_array[634]) begin 
        spike_out_source634 = spike_out_source_array[634];
    end
    always @(spike_out_source_array[635]) begin 
        spike_out_source635 = spike_out_source_array[635];
    end
    always @(spike_out_source_array[636]) begin 
        spike_out_source636 = spike_out_source_array[636];
    end
    always @(spike_out_source_array[637]) begin 
        spike_out_source637 = spike_out_source_array[637];
    end
    always @(spike_out_source_array[638]) begin 
        spike_out_source638 = spike_out_source_array[638];
    end
    always @(spike_out_source_array[639]) begin 
        spike_out_source639 = spike_out_source_array[639];
    end
    always @(spike_out_source_array[640]) begin 
        spike_out_source640 = spike_out_source_array[640];
    end
    always @(spike_out_source_array[641]) begin 
        spike_out_source641 = spike_out_source_array[641];
    end
    always @(spike_out_source_array[642]) begin 
        spike_out_source642 = spike_out_source_array[642];
    end
    always @(spike_out_source_array[643]) begin 
        spike_out_source643 = spike_out_source_array[643];
    end
    always @(spike_out_source_array[644]) begin 
        spike_out_source644 = spike_out_source_array[644];
    end
    always @(spike_out_source_array[645]) begin 
        spike_out_source645 = spike_out_source_array[645];
    end
    always @(spike_out_source_array[646]) begin 
        spike_out_source646 = spike_out_source_array[646];
    end
    always @(spike_out_source_array[647]) begin 
        spike_out_source647 = spike_out_source_array[647];
    end
    always @(spike_out_source_array[648]) begin 
        spike_out_source648 = spike_out_source_array[648];
    end
    always @(spike_out_source_array[649]) begin 
        spike_out_source649 = spike_out_source_array[649];
    end
    always @(spike_out_source_array[650]) begin 
        spike_out_source650 = spike_out_source_array[650];
    end
    always @(spike_out_source_array[651]) begin 
        spike_out_source651 = spike_out_source_array[651];
    end
    always @(spike_out_source_array[652]) begin 
        spike_out_source652 = spike_out_source_array[652];
    end
    always @(spike_out_source_array[653]) begin 
        spike_out_source653 = spike_out_source_array[653];
    end
    always @(spike_out_source_array[654]) begin 
        spike_out_source654 = spike_out_source_array[654];
    end
    always @(spike_out_source_array[655]) begin 
        spike_out_source655 = spike_out_source_array[655];
    end
    always @(spike_out_source_array[656]) begin 
        spike_out_source656 = spike_out_source_array[656];
    end
    always @(spike_out_source_array[657]) begin 
        spike_out_source657 = spike_out_source_array[657];
    end
    always @(spike_out_source_array[658]) begin 
        spike_out_source658 = spike_out_source_array[658];
    end
    always @(spike_out_source_array[659]) begin 
        spike_out_source659 = spike_out_source_array[659];
    end
    always @(spike_out_source_array[660]) begin 
        spike_out_source660 = spike_out_source_array[660];
    end
    always @(spike_out_source_array[661]) begin 
        spike_out_source661 = spike_out_source_array[661];
    end
    always @(spike_out_source_array[662]) begin 
        spike_out_source662 = spike_out_source_array[662];
    end
    always @(spike_out_source_array[663]) begin 
        spike_out_source663 = spike_out_source_array[663];
    end
    always @(spike_out_source_array[664]) begin 
        spike_out_source664 = spike_out_source_array[664];
    end
    always @(spike_out_source_array[665]) begin 
        spike_out_source665 = spike_out_source_array[665];
    end
    always @(spike_out_source_array[666]) begin 
        spike_out_source666 = spike_out_source_array[666];
    end
    always @(spike_out_source_array[667]) begin 
        spike_out_source667 = spike_out_source_array[667];
    end
    always @(spike_out_source_array[668]) begin 
        spike_out_source668 = spike_out_source_array[668];
    end
    always @(spike_out_source_array[669]) begin 
        spike_out_source669 = spike_out_source_array[669];
    end
    always @(spike_out_source_array[670]) begin 
        spike_out_source670 = spike_out_source_array[670];
    end
    always @(spike_out_source_array[671]) begin 
        spike_out_source671 = spike_out_source_array[671];
    end
    always @(spike_out_source_array[672]) begin 
        spike_out_source672 = spike_out_source_array[672];
    end
    always @(spike_out_source_array[673]) begin 
        spike_out_source673 = spike_out_source_array[673];
    end
    always @(spike_out_source_array[674]) begin 
        spike_out_source674 = spike_out_source_array[674];
    end
    always @(spike_out_source_array[675]) begin 
        spike_out_source675 = spike_out_source_array[675];
    end
    always @(spike_out_source_array[676]) begin 
        spike_out_source676 = spike_out_source_array[676];
    end
    always @(spike_out_source_array[677]) begin 
        spike_out_source677 = spike_out_source_array[677];
    end
    always @(spike_out_source_array[678]) begin 
        spike_out_source678 = spike_out_source_array[678];
    end
    always @(spike_out_source_array[679]) begin 
        spike_out_source679 = spike_out_source_array[679];
    end
    always @(spike_out_source_array[680]) begin 
        spike_out_source680 = spike_out_source_array[680];
    end
    always @(spike_out_source_array[681]) begin 
        spike_out_source681 = spike_out_source_array[681];
    end
    always @(spike_out_source_array[682]) begin 
        spike_out_source682 = spike_out_source_array[682];
    end
    always @(spike_out_source_array[683]) begin 
        spike_out_source683 = spike_out_source_array[683];
    end
    always @(spike_out_source_array[684]) begin 
        spike_out_source684 = spike_out_source_array[684];
    end
    always @(spike_out_source_array[685]) begin 
        spike_out_source685 = spike_out_source_array[685];
    end
    always @(spike_out_source_array[686]) begin 
        spike_out_source686 = spike_out_source_array[686];
    end
    always @(spike_out_source_array[687]) begin 
        spike_out_source687 = spike_out_source_array[687];
    end
    always @(spike_out_source_array[688]) begin 
        spike_out_source688 = spike_out_source_array[688];
    end
    always @(spike_out_source_array[689]) begin 
        spike_out_source689 = spike_out_source_array[689];
    end
    always @(spike_out_source_array[690]) begin 
        spike_out_source690 = spike_out_source_array[690];
    end
    always @(spike_out_source_array[691]) begin 
        spike_out_source691 = spike_out_source_array[691];
    end
    always @(spike_out_source_array[692]) begin 
        spike_out_source692 = spike_out_source_array[692];
    end
    always @(spike_out_source_array[693]) begin 
        spike_out_source693 = spike_out_source_array[693];
    end
    always @(spike_out_source_array[694]) begin 
        spike_out_source694 = spike_out_source_array[694];
    end
    always @(spike_out_source_array[695]) begin 
        spike_out_source695 = spike_out_source_array[695];
    end
    always @(spike_out_source_array[696]) begin 
        spike_out_source696 = spike_out_source_array[696];
    end
    always @(spike_out_source_array[697]) begin 
        spike_out_source697 = spike_out_source_array[697];
    end
    always @(spike_out_source_array[698]) begin 
        spike_out_source698 = spike_out_source_array[698];
    end
    always @(spike_out_source_array[699]) begin 
        spike_out_source699 = spike_out_source_array[699];
    end
    always @(spike_out_source_array[700]) begin 
        spike_out_source700 = spike_out_source_array[700];
    end
    always @(spike_out_source_array[701]) begin 
        spike_out_source701 = spike_out_source_array[701];
    end
    always @(spike_out_source_array[702]) begin 
        spike_out_source702 = spike_out_source_array[702];
    end
    always @(spike_out_source_array[703]) begin 
        spike_out_source703 = spike_out_source_array[703];
    end
    always @(spike_out_source_array[704]) begin 
        spike_out_source704 = spike_out_source_array[704];
    end
    always @(spike_out_source_array[705]) begin 
        spike_out_source705 = spike_out_source_array[705];
    end
    always @(spike_out_source_array[706]) begin 
        spike_out_source706 = spike_out_source_array[706];
    end
    always @(spike_out_source_array[707]) begin 
        spike_out_source707 = spike_out_source_array[707];
    end
    always @(spike_out_source_array[708]) begin 
        spike_out_source708 = spike_out_source_array[708];
    end
    always @(spike_out_source_array[709]) begin 
        spike_out_source709 = spike_out_source_array[709];
    end
    always @(spike_out_source_array[710]) begin 
        spike_out_source710 = spike_out_source_array[710];
    end
    always @(spike_out_source_array[711]) begin 
        spike_out_source711 = spike_out_source_array[711];
    end
    always @(spike_out_source_array[712]) begin 
        spike_out_source712 = spike_out_source_array[712];
    end
    always @(spike_out_source_array[713]) begin 
        spike_out_source713 = spike_out_source_array[713];
    end
    always @(spike_out_source_array[714]) begin 
        spike_out_source714 = spike_out_source_array[714];
    end
    always @(spike_out_source_array[715]) begin 
        spike_out_source715 = spike_out_source_array[715];
    end
    always @(spike_out_source_array[716]) begin 
        spike_out_source716 = spike_out_source_array[716];
    end
    always @(spike_out_source_array[717]) begin 
        spike_out_source717 = spike_out_source_array[717];
    end
    always @(spike_out_source_array[718]) begin 
        spike_out_source718 = spike_out_source_array[718];
    end
    always @(spike_out_source_array[719]) begin 
        spike_out_source719 = spike_out_source_array[719];
    end
    always @(spike_out_source_array[720]) begin 
        spike_out_source720 = spike_out_source_array[720];
    end
    always @(spike_out_source_array[721]) begin 
        spike_out_source721 = spike_out_source_array[721];
    end
    always @(spike_out_source_array[722]) begin 
        spike_out_source722 = spike_out_source_array[722];
    end
    always @(spike_out_source_array[723]) begin 
        spike_out_source723 = spike_out_source_array[723];
    end
    always @(spike_out_source_array[724]) begin 
        spike_out_source724 = spike_out_source_array[724];
    end
    always @(spike_out_source_array[725]) begin 
        spike_out_source725 = spike_out_source_array[725];
    end
    always @(spike_out_source_array[726]) begin 
        spike_out_source726 = spike_out_source_array[726];
    end
    always @(spike_out_source_array[727]) begin 
        spike_out_source727 = spike_out_source_array[727];
    end
    always @(spike_out_source_array[728]) begin 
        spike_out_source728 = spike_out_source_array[728];
    end
    always @(spike_out_source_array[729]) begin 
        spike_out_source729 = spike_out_source_array[729];
    end
    always @(spike_out_source_array[730]) begin 
        spike_out_source730 = spike_out_source_array[730];
    end
    always @(spike_out_source_array[731]) begin 
        spike_out_source731 = spike_out_source_array[731];
    end
    always @(spike_out_source_array[732]) begin 
        spike_out_source732 = spike_out_source_array[732];
    end
    always @(spike_out_source_array[733]) begin 
        spike_out_source733 = spike_out_source_array[733];
    end
    always @(spike_out_source_array[734]) begin 
        spike_out_source734 = spike_out_source_array[734];
    end
    always @(spike_out_source_array[735]) begin 
        spike_out_source735 = spike_out_source_array[735];
    end
    always @(spike_out_source_array[736]) begin 
        spike_out_source736 = spike_out_source_array[736];
    end
    always @(spike_out_source_array[737]) begin 
        spike_out_source737 = spike_out_source_array[737];
    end
    always @(spike_out_source_array[738]) begin 
        spike_out_source738 = spike_out_source_array[738];
    end
    always @(spike_out_source_array[739]) begin 
        spike_out_source739 = spike_out_source_array[739];
    end
    always @(spike_out_source_array[740]) begin 
        spike_out_source740 = spike_out_source_array[740];
    end
    always @(spike_out_source_array[741]) begin 
        spike_out_source741 = spike_out_source_array[741];
    end
    always @(spike_out_source_array[742]) begin 
        spike_out_source742 = spike_out_source_array[742];
    end
    always @(spike_out_source_array[743]) begin 
        spike_out_source743 = spike_out_source_array[743];
    end
    always @(spike_out_source_array[744]) begin 
        spike_out_source744 = spike_out_source_array[744];
    end
    always @(spike_out_source_array[745]) begin 
        spike_out_source745 = spike_out_source_array[745];
    end
    always @(spike_out_source_array[746]) begin 
        spike_out_source746 = spike_out_source_array[746];
    end
    always @(spike_out_source_array[747]) begin 
        spike_out_source747 = spike_out_source_array[747];
    end
    always @(spike_out_source_array[748]) begin 
        spike_out_source748 = spike_out_source_array[748];
    end
    always @(spike_out_source_array[749]) begin 
        spike_out_source749 = spike_out_source_array[749];
    end
    always @(spike_out_source_array[750]) begin 
        spike_out_source750 = spike_out_source_array[750];
    end
    always @(spike_out_source_array[751]) begin 
        spike_out_source751 = spike_out_source_array[751];
    end
    always @(spike_out_source_array[752]) begin 
        spike_out_source752 = spike_out_source_array[752];
    end
    always @(spike_out_source_array[753]) begin 
        spike_out_source753 = spike_out_source_array[753];
    end
    always @(spike_out_source_array[754]) begin 
        spike_out_source754 = spike_out_source_array[754];
    end
    always @(spike_out_source_array[755]) begin 
        spike_out_source755 = spike_out_source_array[755];
    end
    always @(spike_out_source_array[756]) begin 
        spike_out_source756 = spike_out_source_array[756];
    end
    always @(spike_out_source_array[757]) begin 
        spike_out_source757 = spike_out_source_array[757];
    end
    always @(spike_out_source_array[758]) begin 
        spike_out_source758 = spike_out_source_array[758];
    end
    always @(spike_out_source_array[759]) begin 
        spike_out_source759 = spike_out_source_array[759];
    end
    always @(spike_out_source_array[760]) begin 
        spike_out_source760 = spike_out_source_array[760];
    end
    always @(spike_out_source_array[761]) begin 
        spike_out_source761 = spike_out_source_array[761];
    end
    always @(spike_out_source_array[762]) begin 
        spike_out_source762 = spike_out_source_array[762];
    end
    always @(spike_out_source_array[763]) begin 
        spike_out_source763 = spike_out_source_array[763];
    end
    always @(spike_out_source_array[764]) begin 
        spike_out_source764 = spike_out_source_array[764];
    end
    always @(spike_out_source_array[765]) begin 
        spike_out_source765 = spike_out_source_array[765];
    end
    always @(spike_out_source_array[766]) begin 
        spike_out_source766 = spike_out_source_array[766];
    end
    always @(spike_out_source_array[767]) begin 
        spike_out_source767 = spike_out_source_array[767];
    end
    always @(spike_out_source_array[768]) begin 
        spike_out_source768 = spike_out_source_array[768];
    end
    always @(spike_out_source_array[769]) begin 
        spike_out_source769 = spike_out_source_array[769];
    end
    always @(spike_out_source_array[770]) begin 
        spike_out_source770 = spike_out_source_array[770];
    end
    always @(spike_out_source_array[771]) begin 
        spike_out_source771 = spike_out_source_array[771];
    end
    always @(spike_out_source_array[772]) begin 
        spike_out_source772 = spike_out_source_array[772];
    end
    always @(spike_out_source_array[773]) begin 
        spike_out_source773 = spike_out_source_array[773];
    end
    always @(spike_out_source_array[774]) begin 
        spike_out_source774 = spike_out_source_array[774];
    end
    always @(spike_out_source_array[775]) begin 
        spike_out_source775 = spike_out_source_array[775];
    end
    always @(spike_out_source_array[776]) begin 
        spike_out_source776 = spike_out_source_array[776];
    end
    always @(spike_out_source_array[777]) begin 
        spike_out_source777 = spike_out_source_array[777];
    end
    always @(spike_out_source_array[778]) begin 
        spike_out_source778 = spike_out_source_array[778];
    end
    always @(spike_out_source_array[779]) begin 
        spike_out_source779 = spike_out_source_array[779];
    end
    always @(spike_out_source_array[780]) begin 
        spike_out_source780 = spike_out_source_array[780];
    end
    always @(spike_out_source_array[781]) begin 
        spike_out_source781 = spike_out_source_array[781];
    end
    always @(spike_out_source_array[782]) begin 
        spike_out_source782 = spike_out_source_array[782];
    end
    always @(spike_out_source_array[783]) begin 
        spike_out_source783 = spike_out_source_array[783];
    end
    always @(spike_out_source_array[784]) begin 
        spike_out_source784 = spike_out_source_array[784];
    end
    always @(spike_out_source_array[785]) begin 
        spike_out_source785 = spike_out_source_array[785];
    end
    always @(spike_out_source_array[786]) begin 
        spike_out_source786 = spike_out_source_array[786];
    end
    always @(spike_out_source_array[787]) begin 
        spike_out_source787 = spike_out_source_array[787];
    end
    always @(spike_out_source_array[788]) begin 
        spike_out_source788 = spike_out_source_array[788];
    end
    always @(spike_out_source_array[789]) begin 
        spike_out_source789 = spike_out_source_array[789];
    end
    always @(spike_out_source_array[790]) begin 
        spike_out_source790 = spike_out_source_array[790];
    end
    always @(spike_out_source_array[791]) begin 
        spike_out_source791 = spike_out_source_array[791];
    end
    always @(spike_out_source_array[792]) begin 
        spike_out_source792 = spike_out_source_array[792];
    end
    always @(spike_out_source_array[793]) begin 
        spike_out_source793 = spike_out_source_array[793];
    end
    always @(spike_out_source_array[794]) begin 
        spike_out_source794 = spike_out_source_array[794];
    end
    always @(spike_out_source_array[795]) begin 
        spike_out_source795 = spike_out_source_array[795];
    end
    always @(spike_out_source_array[796]) begin 
        spike_out_source796 = spike_out_source_array[796];
    end
    always @(spike_out_source_array[797]) begin 
        spike_out_source797 = spike_out_source_array[797];
    end
    always @(spike_out_source_array[798]) begin 
        spike_out_source798 = spike_out_source_array[798];
    end
    always @(spike_out_source_array[799]) begin 
        spike_out_source799 = spike_out_source_array[799];
    end
    always @(spike_out_source_array[800]) begin 
        spike_out_source800 = spike_out_source_array[800];
    end
    always @(spike_out_source_array[801]) begin 
        spike_out_source801 = spike_out_source_array[801];
    end
    always @(spike_out_source_array[802]) begin 
        spike_out_source802 = spike_out_source_array[802];
    end
    always @(spike_out_source_array[803]) begin 
        spike_out_source803 = spike_out_source_array[803];
    end
    always @(spike_out_source_array[804]) begin 
        spike_out_source804 = spike_out_source_array[804];
    end
    always @(spike_out_source_array[805]) begin 
        spike_out_source805 = spike_out_source_array[805];
    end
    always @(spike_out_source_array[806]) begin 
        spike_out_source806 = spike_out_source_array[806];
    end
    always @(spike_out_source_array[807]) begin 
        spike_out_source807 = spike_out_source_array[807];
    end
    always @(spike_out_source_array[808]) begin 
        spike_out_source808 = spike_out_source_array[808];
    end
    always @(spike_out_source_array[809]) begin 
        spike_out_source809 = spike_out_source_array[809];
    end
    always @(spike_out_source_array[810]) begin 
        spike_out_source810 = spike_out_source_array[810];
    end
    always @(spike_out_source_array[811]) begin 
        spike_out_source811 = spike_out_source_array[811];
    end
    always @(spike_out_source_array[812]) begin 
        spike_out_source812 = spike_out_source_array[812];
    end
    always @(spike_out_source_array[813]) begin 
        spike_out_source813 = spike_out_source_array[813];
    end
    always @(spike_out_source_array[814]) begin 
        spike_out_source814 = spike_out_source_array[814];
    end
    always @(spike_out_source_array[815]) begin 
        spike_out_source815 = spike_out_source_array[815];
    end
    always @(spike_out_source_array[816]) begin 
        spike_out_source816 = spike_out_source_array[816];
    end
    always @(spike_out_source_array[817]) begin 
        spike_out_source817 = spike_out_source_array[817];
    end
    always @(spike_out_source_array[818]) begin 
        spike_out_source818 = spike_out_source_array[818];
    end
    always @(spike_out_source_array[819]) begin 
        spike_out_source819 = spike_out_source_array[819];
    end
    always @(spike_out_source_array[820]) begin 
        spike_out_source820 = spike_out_source_array[820];
    end
    always @(spike_out_source_array[821]) begin 
        spike_out_source821 = spike_out_source_array[821];
    end
    always @(spike_out_source_array[822]) begin 
        spike_out_source822 = spike_out_source_array[822];
    end
    always @(spike_out_source_array[823]) begin 
        spike_out_source823 = spike_out_source_array[823];
    end
    always @(spike_out_source_array[824]) begin 
        spike_out_source824 = spike_out_source_array[824];
    end
    always @(spike_out_source_array[825]) begin 
        spike_out_source825 = spike_out_source_array[825];
    end
    always @(spike_out_source_array[826]) begin 
        spike_out_source826 = spike_out_source_array[826];
    end
    always @(spike_out_source_array[827]) begin 
        spike_out_source827 = spike_out_source_array[827];
    end
    always @(spike_out_source_array[828]) begin 
        spike_out_source828 = spike_out_source_array[828];
    end
    always @(spike_out_source_array[829]) begin 
        spike_out_source829 = spike_out_source_array[829];
    end
    always @(spike_out_source_array[830]) begin 
        spike_out_source830 = spike_out_source_array[830];
    end
    always @(spike_out_source_array[831]) begin 
        spike_out_source831 = spike_out_source_array[831];
    end
    always @(spike_out_source_array[832]) begin 
        spike_out_source832 = spike_out_source_array[832];
    end
    always @(spike_out_source_array[833]) begin 
        spike_out_source833 = spike_out_source_array[833];
    end
    always @(spike_out_source_array[834]) begin 
        spike_out_source834 = spike_out_source_array[834];
    end
    always @(spike_out_source_array[835]) begin 
        spike_out_source835 = spike_out_source_array[835];
    end
    always @(spike_out_source_array[836]) begin 
        spike_out_source836 = spike_out_source_array[836];
    end
    always @(spike_out_source_array[837]) begin 
        spike_out_source837 = spike_out_source_array[837];
    end
    always @(spike_out_source_array[838]) begin 
        spike_out_source838 = spike_out_source_array[838];
    end
    always @(spike_out_source_array[839]) begin 
        spike_out_source839 = spike_out_source_array[839];
    end
    always @(spike_out_source_array[840]) begin 
        spike_out_source840 = spike_out_source_array[840];
    end
    always @(spike_out_source_array[841]) begin 
        spike_out_source841 = spike_out_source_array[841];
    end
    always @(spike_out_source_array[842]) begin 
        spike_out_source842 = spike_out_source_array[842];
    end
    always @(spike_out_source_array[843]) begin 
        spike_out_source843 = spike_out_source_array[843];
    end
    always @(spike_out_source_array[844]) begin 
        spike_out_source844 = spike_out_source_array[844];
    end
    always @(spike_out_source_array[845]) begin 
        spike_out_source845 = spike_out_source_array[845];
    end
    always @(spike_out_source_array[846]) begin 
        spike_out_source846 = spike_out_source_array[846];
    end
    always @(spike_out_source_array[847]) begin 
        spike_out_source847 = spike_out_source_array[847];
    end
    always @(spike_out_source_array[848]) begin 
        spike_out_source848 = spike_out_source_array[848];
    end
    always @(spike_out_source_array[849]) begin 
        spike_out_source849 = spike_out_source_array[849];
    end
    always @(spike_out_source_array[850]) begin 
        spike_out_source850 = spike_out_source_array[850];
    end
    always @(spike_out_source_array[851]) begin 
        spike_out_source851 = spike_out_source_array[851];
    end
    always @(spike_out_source_array[852]) begin 
        spike_out_source852 = spike_out_source_array[852];
    end
    always @(spike_out_source_array[853]) begin 
        spike_out_source853 = spike_out_source_array[853];
    end
    always @(spike_out_source_array[854]) begin 
        spike_out_source854 = spike_out_source_array[854];
    end
    always @(spike_out_source_array[855]) begin 
        spike_out_source855 = spike_out_source_array[855];
    end
    always @(spike_out_source_array[856]) begin 
        spike_out_source856 = spike_out_source_array[856];
    end
    always @(spike_out_source_array[857]) begin 
        spike_out_source857 = spike_out_source_array[857];
    end
    always @(spike_out_source_array[858]) begin 
        spike_out_source858 = spike_out_source_array[858];
    end
    always @(spike_out_source_array[859]) begin 
        spike_out_source859 = spike_out_source_array[859];
    end
    always @(spike_out_source_array[860]) begin 
        spike_out_source860 = spike_out_source_array[860];
    end
    always @(spike_out_source_array[861]) begin 
        spike_out_source861 = spike_out_source_array[861];
    end
    always @(spike_out_source_array[862]) begin 
        spike_out_source862 = spike_out_source_array[862];
    end
    always @(spike_out_source_array[863]) begin 
        spike_out_source863 = spike_out_source_array[863];
    end
    always @(spike_out_source_array[864]) begin 
        spike_out_source864 = spike_out_source_array[864];
    end
    always @(spike_out_source_array[865]) begin 
        spike_out_source865 = spike_out_source_array[865];
    end
    always @(spike_out_source_array[866]) begin 
        spike_out_source866 = spike_out_source_array[866];
    end
    always @(spike_out_source_array[867]) begin 
        spike_out_source867 = spike_out_source_array[867];
    end
    always @(spike_out_source_array[868]) begin 
        spike_out_source868 = spike_out_source_array[868];
    end
    always @(spike_out_source_array[869]) begin 
        spike_out_source869 = spike_out_source_array[869];
    end
    always @(spike_out_source_array[870]) begin 
        spike_out_source870 = spike_out_source_array[870];
    end
    always @(spike_out_source_array[871]) begin 
        spike_out_source871 = spike_out_source_array[871];
    end
    always @(spike_out_source_array[872]) begin 
        spike_out_source872 = spike_out_source_array[872];
    end
    always @(spike_out_source_array[873]) begin 
        spike_out_source873 = spike_out_source_array[873];
    end
    always @(spike_out_source_array[874]) begin 
        spike_out_source874 = spike_out_source_array[874];
    end
    always @(spike_out_source_array[875]) begin 
        spike_out_source875 = spike_out_source_array[875];
    end
    always @(spike_out_source_array[876]) begin 
        spike_out_source876 = spike_out_source_array[876];
    end
    always @(spike_out_source_array[877]) begin 
        spike_out_source877 = spike_out_source_array[877];
    end
    always @(spike_out_source_array[878]) begin 
        spike_out_source878 = spike_out_source_array[878];
    end
    always @(spike_out_source_array[879]) begin 
        spike_out_source879 = spike_out_source_array[879];
    end
    always @(spike_out_source_array[880]) begin 
        spike_out_source880 = spike_out_source_array[880];
    end
    always @(spike_out_source_array[881]) begin 
        spike_out_source881 = spike_out_source_array[881];
    end
    always @(spike_out_source_array[882]) begin 
        spike_out_source882 = spike_out_source_array[882];
    end
    always @(spike_out_source_array[883]) begin 
        spike_out_source883 = spike_out_source_array[883];
    end
    always @(spike_out_source_array[884]) begin 
        spike_out_source884 = spike_out_source_array[884];
    end
    always @(spike_out_source_array[885]) begin 
        spike_out_source885 = spike_out_source_array[885];
    end
    always @(spike_out_source_array[886]) begin 
        spike_out_source886 = spike_out_source_array[886];
    end
    always @(spike_out_source_array[887]) begin 
        spike_out_source887 = spike_out_source_array[887];
    end
    always @(spike_out_source_array[888]) begin 
        spike_out_source888 = spike_out_source_array[888];
    end
    always @(spike_out_source_array[889]) begin 
        spike_out_source889 = spike_out_source_array[889];
    end
    always @(spike_out_source_array[890]) begin 
        spike_out_source890 = spike_out_source_array[890];
    end
    always @(spike_out_source_array[891]) begin 
        spike_out_source891 = spike_out_source_array[891];
    end
    always @(spike_out_source_array[892]) begin 
        spike_out_source892 = spike_out_source_array[892];
    end
    always @(spike_out_source_array[893]) begin 
        spike_out_source893 = spike_out_source_array[893];
    end
    always @(spike_out_source_array[894]) begin 
        spike_out_source894 = spike_out_source_array[894];
    end
    always @(spike_out_source_array[895]) begin 
        spike_out_source895 = spike_out_source_array[895];
    end
    always @(spike_out_source_array[896]) begin 
        spike_out_source896 = spike_out_source_array[896];
    end
    always @(spike_out_source_array[897]) begin 
        spike_out_source897 = spike_out_source_array[897];
    end
    always @(spike_out_source_array[898]) begin 
        spike_out_source898 = spike_out_source_array[898];
    end
    always @(spike_out_source_array[899]) begin 
        spike_out_source899 = spike_out_source_array[899];
    end
    always @(spike_out_source_array[900]) begin 
        spike_out_source900 = spike_out_source_array[900];
    end
    always @(spike_out_source_array[901]) begin 
        spike_out_source901 = spike_out_source_array[901];
    end
    always @(spike_out_source_array[902]) begin 
        spike_out_source902 = spike_out_source_array[902];
    end
    always @(spike_out_source_array[903]) begin 
        spike_out_source903 = spike_out_source_array[903];
    end
    always @(spike_out_source_array[904]) begin 
        spike_out_source904 = spike_out_source_array[904];
    end
    always @(spike_out_source_array[905]) begin 
        spike_out_source905 = spike_out_source_array[905];
    end
    always @(spike_out_source_array[906]) begin 
        spike_out_source906 = spike_out_source_array[906];
    end
    always @(spike_out_source_array[907]) begin 
        spike_out_source907 = spike_out_source_array[907];
    end
    always @(spike_out_source_array[908]) begin 
        spike_out_source908 = spike_out_source_array[908];
    end
    always @(spike_out_source_array[909]) begin 
        spike_out_source909 = spike_out_source_array[909];
    end
    always @(spike_out_source_array[910]) begin 
        spike_out_source910 = spike_out_source_array[910];
    end
    always @(spike_out_source_array[911]) begin 
        spike_out_source911 = spike_out_source_array[911];
    end
    always @(spike_out_source_array[912]) begin 
        spike_out_source912 = spike_out_source_array[912];
    end
    always @(spike_out_source_array[913]) begin 
        spike_out_source913 = spike_out_source_array[913];
    end
    always @(spike_out_source_array[914]) begin 
        spike_out_source914 = spike_out_source_array[914];
    end
    always @(spike_out_source_array[915]) begin 
        spike_out_source915 = spike_out_source_array[915];
    end
    always @(spike_out_source_array[916]) begin 
        spike_out_source916 = spike_out_source_array[916];
    end
    always @(spike_out_source_array[917]) begin 
        spike_out_source917 = spike_out_source_array[917];
    end
    always @(spike_out_source_array[918]) begin 
        spike_out_source918 = spike_out_source_array[918];
    end
    always @(spike_out_source_array[919]) begin 
        spike_out_source919 = spike_out_source_array[919];
    end
    always @(spike_out_source_array[920]) begin 
        spike_out_source920 = spike_out_source_array[920];
    end
    always @(spike_out_source_array[921]) begin 
        spike_out_source921 = spike_out_source_array[921];
    end
    always @(spike_out_source_array[922]) begin 
        spike_out_source922 = spike_out_source_array[922];
    end
    always @(spike_out_source_array[923]) begin 
        spike_out_source923 = spike_out_source_array[923];
    end
    always @(spike_out_source_array[924]) begin 
        spike_out_source924 = spike_out_source_array[924];
    end
    always @(spike_out_source_array[925]) begin 
        spike_out_source925 = spike_out_source_array[925];
    end
    always @(spike_out_source_array[926]) begin 
        spike_out_source926 = spike_out_source_array[926];
    end
    always @(spike_out_source_array[927]) begin 
        spike_out_source927 = spike_out_source_array[927];
    end
    always @(spike_out_source_array[928]) begin 
        spike_out_source928 = spike_out_source_array[928];
    end
    always @(spike_out_source_array[929]) begin 
        spike_out_source929 = spike_out_source_array[929];
    end
    always @(spike_out_source_array[930]) begin 
        spike_out_source930 = spike_out_source_array[930];
    end
    always @(spike_out_source_array[931]) begin 
        spike_out_source931 = spike_out_source_array[931];
    end
    always @(spike_out_source_array[932]) begin 
        spike_out_source932 = spike_out_source_array[932];
    end
    always @(spike_out_source_array[933]) begin 
        spike_out_source933 = spike_out_source_array[933];
    end
    always @(spike_out_source_array[934]) begin 
        spike_out_source934 = spike_out_source_array[934];
    end
    always @(spike_out_source_array[935]) begin 
        spike_out_source935 = spike_out_source_array[935];
    end
    always @(spike_out_source_array[936]) begin 
        spike_out_source936 = spike_out_source_array[936];
    end
    always @(spike_out_source_array[937]) begin 
        spike_out_source937 = spike_out_source_array[937];
    end
    always @(spike_out_source_array[938]) begin 
        spike_out_source938 = spike_out_source_array[938];
    end
    always @(spike_out_source_array[939]) begin 
        spike_out_source939 = spike_out_source_array[939];
    end
    always @(spike_out_source_array[940]) begin 
        spike_out_source940 = spike_out_source_array[940];
    end
    always @(spike_out_source_array[941]) begin 
        spike_out_source941 = spike_out_source_array[941];
    end
    always @(spike_out_source_array[942]) begin 
        spike_out_source942 = spike_out_source_array[942];
    end
    always @(spike_out_source_array[943]) begin 
        spike_out_source943 = spike_out_source_array[943];
    end
    always @(spike_out_source_array[944]) begin 
        spike_out_source944 = spike_out_source_array[944];
    end
    always @(spike_out_source_array[945]) begin 
        spike_out_source945 = spike_out_source_array[945];
    end
    always @(spike_out_source_array[946]) begin 
        spike_out_source946 = spike_out_source_array[946];
    end
    always @(spike_out_source_array[947]) begin 
        spike_out_source947 = spike_out_source_array[947];
    end
    always @(spike_out_source_array[948]) begin 
        spike_out_source948 = spike_out_source_array[948];
    end
    always @(spike_out_source_array[949]) begin 
        spike_out_source949 = spike_out_source_array[949];
    end
    always @(spike_out_source_array[950]) begin 
        spike_out_source950 = spike_out_source_array[950];
    end
    always @(spike_out_source_array[951]) begin 
        spike_out_source951 = spike_out_source_array[951];
    end
    always @(spike_out_source_array[952]) begin 
        spike_out_source952 = spike_out_source_array[952];
    end
    always @(spike_out_source_array[953]) begin 
        spike_out_source953 = spike_out_source_array[953];
    end
    always @(spike_out_source_array[954]) begin 
        spike_out_source954 = spike_out_source_array[954];
    end
    always @(spike_out_source_array[955]) begin 
        spike_out_source955 = spike_out_source_array[955];
    end
    always @(spike_out_source_array[956]) begin 
        spike_out_source956 = spike_out_source_array[956];
    end
    always @(spike_out_source_array[957]) begin 
        spike_out_source957 = spike_out_source_array[957];
    end
    always @(spike_out_source_array[958]) begin 
        spike_out_source958 = spike_out_source_array[958];
    end
    always @(spike_out_source_array[959]) begin 
        spike_out_source959 = spike_out_source_array[959];
    end
    always @(spike_out_source_array[960]) begin 
        spike_out_source960 = spike_out_source_array[960];
    end
    always @(spike_out_source_array[961]) begin 
        spike_out_source961 = spike_out_source_array[961];
    end
    always @(spike_out_source_array[962]) begin 
        spike_out_source962 = spike_out_source_array[962];
    end
    always @(spike_out_source_array[963]) begin 
        spike_out_source963 = spike_out_source_array[963];
    end
    always @(spike_out_source_array[964]) begin 
        spike_out_source964 = spike_out_source_array[964];
    end
    always @(spike_out_source_array[965]) begin 
        spike_out_source965 = spike_out_source_array[965];
    end
    always @(spike_out_source_array[966]) begin 
        spike_out_source966 = spike_out_source_array[966];
    end
    always @(spike_out_source_array[967]) begin 
        spike_out_source967 = spike_out_source_array[967];
    end
    always @(spike_out_source_array[968]) begin 
        spike_out_source968 = spike_out_source_array[968];
    end
    always @(spike_out_source_array[969]) begin 
        spike_out_source969 = spike_out_source_array[969];
    end
    always @(spike_out_source_array[970]) begin 
        spike_out_source970 = spike_out_source_array[970];
    end
    always @(spike_out_source_array[971]) begin 
        spike_out_source971 = spike_out_source_array[971];
    end
    always @(spike_out_source_array[972]) begin 
        spike_out_source972 = spike_out_source_array[972];
    end
    always @(spike_out_source_array[973]) begin 
        spike_out_source973 = spike_out_source_array[973];
    end
    always @(spike_out_source_array[974]) begin 
        spike_out_source974 = spike_out_source_array[974];
    end
    always @(spike_out_source_array[975]) begin 
        spike_out_source975 = spike_out_source_array[975];
    end
    always @(spike_out_source_array[976]) begin 
        spike_out_source976 = spike_out_source_array[976];
    end
    always @(spike_out_source_array[977]) begin 
        spike_out_source977 = spike_out_source_array[977];
    end
    always @(spike_out_source_array[978]) begin 
        spike_out_source978 = spike_out_source_array[978];
    end
    always @(spike_out_source_array[979]) begin 
        spike_out_source979 = spike_out_source_array[979];
    end
    always @(spike_out_source_array[980]) begin 
        spike_out_source980 = spike_out_source_array[980];
    end
    always @(spike_out_source_array[981]) begin 
        spike_out_source981 = spike_out_source_array[981];
    end
    always @(spike_out_source_array[982]) begin 
        spike_out_source982 = spike_out_source_array[982];
    end
    always @(spike_out_source_array[983]) begin 
        spike_out_source983 = spike_out_source_array[983];
    end
    always @(spike_out_source_array[984]) begin 
        spike_out_source984 = spike_out_source_array[984];
    end
    always @(spike_out_source_array[985]) begin 
        spike_out_source985 = spike_out_source_array[985];
    end
    always @(spike_out_source_array[986]) begin 
        spike_out_source986 = spike_out_source_array[986];
    end
    always @(spike_out_source_array[987]) begin 
        spike_out_source987 = spike_out_source_array[987];
    end
    always @(spike_out_source_array[988]) begin 
        spike_out_source988 = spike_out_source_array[988];
    end
    always @(spike_out_source_array[989]) begin 
        spike_out_source989 = spike_out_source_array[989];
    end
    always @(spike_out_source_array[990]) begin 
        spike_out_source990 = spike_out_source_array[990];
    end
    always @(spike_out_source_array[991]) begin 
        spike_out_source991 = spike_out_source_array[991];
    end
    always @(spike_out_source_array[992]) begin 
        spike_out_source992 = spike_out_source_array[992];
    end
    always @(spike_out_source_array[993]) begin 
        spike_out_source993 = spike_out_source_array[993];
    end
    always @(spike_out_source_array[994]) begin 
        spike_out_source994 = spike_out_source_array[994];
    end
    always @(spike_out_source_array[995]) begin 
        spike_out_source995 = spike_out_source_array[995];
    end
    always @(spike_out_source_array[996]) begin 
        spike_out_source996 = spike_out_source_array[996];
    end
    always @(spike_out_source_array[997]) begin 
        spike_out_source997 = spike_out_source_array[997];
    end
    always @(spike_out_source_array[998]) begin 
        spike_out_source998 = spike_out_source_array[998];
    end
    always @(spike_out_source_array[999]) begin 
        spike_out_source999 = spike_out_source_array[999];
    end
    always @(spike_out_source_array[1000]) begin 
        spike_out_source1000 = spike_out_source_array[1000];
    end
    always @(spike_out_source_array[1001]) begin 
        spike_out_source1001 = spike_out_source_array[1001];
    end
    always @(spike_out_source_array[1002]) begin 
        spike_out_source1002 = spike_out_source_array[1002];
    end
    always @(spike_out_source_array[1003]) begin 
        spike_out_source1003 = spike_out_source_array[1003];
    end
    always @(spike_out_source_array[1004]) begin 
        spike_out_source1004 = spike_out_source_array[1004];
    end
    always @(spike_out_source_array[1005]) begin 
        spike_out_source1005 = spike_out_source_array[1005];
    end
    always @(spike_out_source_array[1006]) begin 
        spike_out_source1006 = spike_out_source_array[1006];
    end
    always @(spike_out_source_array[1007]) begin 
        spike_out_source1007 = spike_out_source_array[1007];
    end
    always @(spike_out_source_array[1008]) begin 
        spike_out_source1008 = spike_out_source_array[1008];
    end
    always @(spike_out_source_array[1009]) begin 
        spike_out_source1009 = spike_out_source_array[1009];
    end
    always @(spike_out_source_array[1010]) begin 
        spike_out_source1010 = spike_out_source_array[1010];
    end
    always @(spike_out_source_array[1011]) begin 
        spike_out_source1011 = spike_out_source_array[1011];
    end
    always @(spike_out_source_array[1012]) begin 
        spike_out_source1012 = spike_out_source_array[1012];
    end
    always @(spike_out_source_array[1013]) begin 
        spike_out_source1013 = spike_out_source_array[1013];
    end
    always @(spike_out_source_array[1014]) begin 
        spike_out_source1014 = spike_out_source_array[1014];
    end
    always @(spike_out_source_array[1015]) begin 
        spike_out_source1015 = spike_out_source_array[1015];
    end
    always @(spike_out_source_array[1016]) begin 
        spike_out_source1016 = spike_out_source_array[1016];
    end
    always @(spike_out_source_array[1017]) begin 
        spike_out_source1017 = spike_out_source_array[1017];
    end
    always @(spike_out_source_array[1018]) begin 
        spike_out_source1018 = spike_out_source_array[1018];
    end
    always @(spike_out_source_array[1019]) begin 
        spike_out_source1019 = spike_out_source_array[1019];
    end
    always @(spike_out_source_array[1020]) begin 
        spike_out_source1020 = spike_out_source_array[1020];
    end
    always @(spike_out_source_array[1021]) begin 
        spike_out_source1021 = spike_out_source_array[1021];
    end
    always @(spike_out_source_array[1022]) begin 
        spike_out_source1022 = spike_out_source_array[1022];
    end
    always @(spike_out_source_array[1023]) begin 
        spike_out_source1023 = spike_out_source_array[1023];
    end
    reg[18:0] i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21, module network_interface_scaled (
        input wire spike0,
    input wire spike1,    input wire spike2,    input wire spike3,    input wire spike4,    input wire spike5,    input wire spike6,    input wire spike7,    input wire spike8,    input wire spike9,    input wire spike10,    input wire spike11,    input wire spike12,    input wire spike13,    input wire spike14,    input wire spike15,    input wire spike16,    input wire spike17,    input wire spike18,    input wire spike19,    input wire spike20,    input wire spike21,    input wire spike22,    input wire spike23,    input wire spike24,    input wire spike25,    input wire spike26,    input wire spike27,    input wire spike28,    input wire spike29,    input wire spike30,    input wire spike31,    input wire spike32,    input wire spike33,    input wire spike34,    input wire spike35,    input wire spike36,    input wire spike37,    input wire spike38,    input wire spike39,    input wire spike40,    input wire spike41,    input wire spike42,    input wire spike43,    input wire spike44,    input wire spike45,    input wire spike46,    input wire spike47,    input wire spike48,    input wire spike49,    input wire spike50,    input wire spike51,    input wire spike52,    input wire spike53,    input wire spike54,    input wire spike55,    input wire spike56,    input wire spike57,    input wire spike58,    input wire spike59,    input wire spike60,    input wire spike61,    input wire spike62,    input wire spike63,    input wire spike64,    input wire spike65,    input wire spike66,    input wire spike67,    input wire spike68,    input wire spike69,    input wire spike70,    input wire spike71,    input wire spike72,    input wire spike73,    input wire spike74,    input wire spike75,    input wire spike76,    input wire spike77,    input wire spike78,    input wire spike79,    input wire spike80,    input wire spike81,    input wire spike82,    input wire spike83,    input wire spike84,    input wire spike85,    input wire spike86,    input wire spike87,    input wire spike88,    input wire spike89,    input wire spike90,    input wire spike91,    input wire spike92,    input wire spike93,    input wire spike94,    input wire spike95,    input wire spike96,    input wire spike97,    input wire spike98,    input wire spike99,    input wire spike100,
    input wire spike101,    input wire spike102,    input wire spike103,    input wire spike104,    input wire spike105,    input wire spike106,    input wire spike107,    input wire spike108,    input wire spike109,    input wire spike110,    input wire spike111,    input wire spike112,    input wire spike113,    input wire spike114,    input wire spike115,    input wire spike116,    input wire spike117,    input wire spike118,    input wire spike119,    input wire spike120,    input wire spike121,    input wire spike122,    input wire spike123,    input wire spike124,    input wire spike125,    input wire spike126,    input wire spike127,    input wire spike128,    input wire spike129,    input wire spike130,    input wire spike131,    input wire spike132,    input wire spike133,    input wire spike134,    input wire spike135,    input wire spike136,    input wire spike137,    input wire spike138,    input wire spike139,    input wire spike140,    input wire spike141,    input wire spike142,    input wire spike143,    input wire spike144,    input wire spike145,    input wire spike146,    input wire spike147,    input wire spike148,    input wire spike149,    input wire spike150,    input wire spike151,    input wire spike152,    input wire spike153,    input wire spike154,    input wire spike155,    input wire spike156,    input wire spike157,    input wire spike158,    input wire spike159,    input wire spike160,    input wire spike161,    input wire spike162,    input wire spike163,    input wire spike164,    input wire spike165,    input wire spike166,    input wire spike167,    input wire spike168,    input wire spike169,    input wire spike170,    input wire spike171,    input wire spike172,    input wire spike173,    input wire spike174,    input wire spike175,    input wire spike176,    input wire spike177,    input wire spike178,    input wire spike179,    input wire spike180,    input wire spike181,    input wire spike182,    input wire spike183,    input wire spike184,    input wire spike185,    input wire spike186,    input wire spike187,    input wire spike188,    input wire spike189,    input wire spike190,    input wire spike191,    input wire spike192,    input wire spike193,    input wire spike194,    input wire spike195,    input wire spike196,    input wire spike197,    input wire spike198,    input wire spike199,    input wire spike200,
    input wire spike201,    input wire spike202,    input wire spike203,    input wire spike204,    input wire spike205,    input wire spike206,    input wire spike207,    input wire spike208,    input wire spike209,    input wire spike210,    input wire spike211,    input wire spike212,    input wire spike213,    input wire spike214,    input wire spike215,    input wire spike216,    input wire spike217,    input wire spike218,    input wire spike219,    input wire spike220,    input wire spike221,    input wire spike222,    input wire spike223,    input wire spike224,    input wire spike225,    input wire spike226,    input wire spike227,    input wire spike228,    input wire spike229,    input wire spike230,    input wire spike231,    input wire spike232,    input wire spike233,    input wire spike234,    input wire spike235,    input wire spike236,    input wire spike237,    input wire spike238,    input wire spike239,    input wire spike240,    input wire spike241,    input wire spike242,    input wire spike243,    input wire spike244,    input wire spike245,    input wire spike246,    input wire spike247,    input wire spike248,    input wire spike249,    input wire spike250,    input wire spike251,    input wire spike252,    input wire spike253,    input wire spike254,    input wire spike255,    input wire spike256,    input wire spike257,    input wire spike258,    input wire spike259,    input wire spike260,    input wire spike261,    input wire spike262,    input wire spike263,    input wire spike264,    input wire spike265,    input wire spike266,    input wire spike267,    input wire spike268,    input wire spike269,    input wire spike270,    input wire spike271,    input wire spike272,    input wire spike273,    input wire spike274,    input wire spike275,    input wire spike276,    input wire spike277,    input wire spike278,    input wire spike279,    input wire spike280,    input wire spike281,    input wire spike282,    input wire spike283,    input wire spike284,    input wire spike285,    input wire spike286,    input wire spike287,    input wire spike288,    input wire spike289,    input wire spike290,    input wire spike291,    input wire spike292,    input wire spike293,    input wire spike294,    input wire spike295,    input wire spike296,    input wire spike297,    input wire spike298,    input wire spike299,    input wire spike300,
    input wire spike301,    input wire spike302,    input wire spike303,    input wire spike304,    input wire spike305,    input wire spike306,    input wire spike307,    input wire spike308,    input wire spike309,    input wire spike310,    input wire spike311,    input wire spike312,    input wire spike313,    input wire spike314,    input wire spike315,    input wire spike316,    input wire spike317,    input wire spike318,    input wire spike319,    input wire spike320,    input wire spike321,    input wire spike322,    input wire spike323,    input wire spike324,    input wire spike325,    input wire spike326,    input wire spike327,    input wire spike328,    input wire spike329,    input wire spike330,    input wire spike331,    input wire spike332,    input wire spike333,    input wire spike334,    input wire spike335,    input wire spike336,    input wire spike337,    input wire spike338,    input wire spike339,    input wire spike340,    input wire spike341,    input wire spike342,    input wire spike343,    input wire spike344,    input wire spike345,    input wire spike346,    input wire spike347,    input wire spike348,    input wire spike349,    input wire spike350,    input wire spike351,    input wire spike352,    input wire spike353,    input wire spike354,    input wire spike355,    input wire spike356,    input wire spike357,    input wire spike358,    input wire spike359,    input wire spike360,    input wire spike361,    input wire spike362,    input wire spike363,    input wire spike364,    input wire spike365,    input wire spike366,    input wire spike367,    input wire spike368,    input wire spike369,    input wire spike370,    input wire spike371,    input wire spike372,    input wire spike373,    input wire spike374,    input wire spike375,    input wire spike376,    input wire spike377,    input wire spike378,    input wire spike379,    input wire spike380,    input wire spike381,    input wire spike382,    input wire spike383,    input wire spike384,    input wire spike385,    input wire spike386,    input wire spike387,    input wire spike388,    input wire spike389,    input wire spike390,    input wire spike391,    input wire spike392,    input wire spike393,    input wire spike394,    input wire spike395,    input wire spike396,    input wire spike397,    input wire spike398,    input wire spike399,    input wire spike400,
    input wire spike401,    input wire spike402,    input wire spike403,    input wire spike404,    input wire spike405,    input wire spike406,    input wire spike407,    input wire spike408,    input wire spike409,    input wire spike410,    input wire spike411,    input wire spike412,    input wire spike413,    input wire spike414,    input wire spike415,    input wire spike416,    input wire spike417,    input wire spike418,    input wire spike419,    input wire spike420,    input wire spike421,    input wire spike422,    input wire spike423,    input wire spike424,    input wire spike425,    input wire spike426,    input wire spike427,    input wire spike428,    input wire spike429,    input wire spike430,    input wire spike431,    input wire spike432,    input wire spike433,    input wire spike434,    input wire spike435,    input wire spike436,    input wire spike437,    input wire spike438,    input wire spike439,    input wire spike440,    input wire spike441,    input wire spike442,    input wire spike443,    input wire spike444,    input wire spike445,    input wire spike446,    input wire spike447,    input wire spike448,    input wire spike449,    input wire spike450,    input wire spike451,    input wire spike452,    input wire spike453,    input wire spike454,    input wire spike455,    input wire spike456,    input wire spike457,    input wire spike458,    input wire spike459,    input wire spike460,    input wire spike461,    input wire spike462,    input wire spike463,    input wire spike464,    input wire spike465,    input wire spike466,    input wire spike467,    input wire spike468,    input wire spike469,    input wire spike470,    input wire spike471,    input wire spike472,    input wire spike473,    input wire spike474,    input wire spike475,    input wire spike476,    input wire spike477,    input wire spike478,    input wire spike479,    input wire spike480,    input wire spike481,    input wire spike482,    input wire spike483,    input wire spike484,    input wire spike485,    input wire spike486,    input wire spike487,    input wire spike488,    input wire spike489,    input wire spike490,    input wire spike491,    input wire spike492,    input wire spike493,    input wire spike494,    input wire spike495,    input wire spike496,    input wire spike497,    input wire spike498,    input wire spike499,    input wire spike500,
    input wire spike501,    input wire spike502,    input wire spike503,    input wire spike504,    input wire spike505,    input wire spike506,    input wire spike507,    input wire spike508,    input wire spike509,    input wire spike510,    input wire spike511,    input wire spike512,    input wire spike513,    input wire spike514,    input wire spike515,    input wire spike516,    input wire spike517,    input wire spike518,    input wire spike519,    input wire spike520,    input wire spike521,    input wire spike522,    input wire spike523,    input wire spike524,    input wire spike525,    input wire spike526,    input wire spike527,    input wire spike528,    input wire spike529,    input wire spike530,    input wire spike531,    input wire spike532,    input wire spike533,    input wire spike534,    input wire spike535,    input wire spike536,    input wire spike537,    input wire spike538,    input wire spike539,    input wire spike540,    input wire spike541,    input wire spike542,    input wire spike543,    input wire spike544,    input wire spike545,    input wire spike546,    input wire spike547,    input wire spike548,    input wire spike549,    input wire spike550,    input wire spike551,    input wire spike552,    input wire spike553,    input wire spike554,    input wire spike555,    input wire spike556,    input wire spike557,    input wire spike558,    input wire spike559,    input wire spike560,    input wire spike561,    input wire spike562,    input wire spike563,    input wire spike564,    input wire spike565,    input wire spike566,    input wire spike567,    input wire spike568,    input wire spike569,    input wire spike570,    input wire spike571,    input wire spike572,    input wire spike573,    input wire spike574,    input wire spike575,    input wire spike576,    input wire spike577,    input wire spike578,    input wire spike579,    input wire spike580,    input wire spike581,    input wire spike582,    input wire spike583,    input wire spike584,    input wire spike585,    input wire spike586,    input wire spike587,    input wire spike588,    input wire spike589,    input wire spike590,    input wire spike591,    input wire spike592,    input wire spike593,    input wire spike594,    input wire spike595,    input wire spike596,    input wire spike597,    input wire spike598,    input wire spike599,    input wire spike600,
    input wire spike601,    input wire spike602,    input wire spike603,    input wire spike604,    input wire spike605,    input wire spike606,    input wire spike607,    input wire spike608,    input wire spike609,    input wire spike610,    input wire spike611,    input wire spike612,    input wire spike613,    input wire spike614,    input wire spike615,    input wire spike616,    input wire spike617,    input wire spike618,    input wire spike619,    input wire spike620,    input wire spike621,    input wire spike622,    input wire spike623,    input wire spike624,    input wire spike625,    input wire spike626,    input wire spike627,    input wire spike628,    input wire spike629,    input wire spike630,    input wire spike631,    input wire spike632,    input wire spike633,    input wire spike634,    input wire spike635,    input wire spike636,    input wire spike637,    input wire spike638,    input wire spike639,    input wire spike640,    input wire spike641,    input wire spike642,    input wire spike643,    input wire spike644,    input wire spike645,    input wire spike646,    input wire spike647,    input wire spike648,    input wire spike649,    input wire spike650,    input wire spike651,    input wire spike652,    input wire spike653,    input wire spike654,    input wire spike655,    input wire spike656,    input wire spike657,    input wire spike658,    input wire spike659,    input wire spike660,    input wire spike661,    input wire spike662,    input wire spike663,    input wire spike664,    input wire spike665,    input wire spike666,    input wire spike667,    input wire spike668,    input wire spike669,    input wire spike670,    input wire spike671,    input wire spike672,    input wire spike673,    input wire spike674,    input wire spike675,    input wire spike676,    input wire spike677,    input wire spike678,    input wire spike679,    input wire spike680,    input wire spike681,    input wire spike682,    input wire spike683,    input wire spike684,    input wire spike685,    input wire spike686,    input wire spike687,    input wire spike688,    input wire spike689,    input wire spike690,    input wire spike691,    input wire spike692,    input wire spike693,    input wire spike694,    input wire spike695,    input wire spike696,    input wire spike697,    input wire spike698,    input wire spike699,    input wire spike700,
    input wire spike701,    input wire spike702,    input wire spike703,    input wire spike704,    input wire spike705,    input wire spike706,    input wire spike707,    input wire spike708,    input wire spike709,    input wire spike710,    input wire spike711,    input wire spike712,    input wire spike713,    input wire spike714,    input wire spike715,    input wire spike716,    input wire spike717,    input wire spike718,    input wire spike719,    input wire spike720,    input wire spike721,    input wire spike722,    input wire spike723,    input wire spike724,    input wire spike725,    input wire spike726,    input wire spike727,    input wire spike728,    input wire spike729,    input wire spike730,    input wire spike731,    input wire spike732,    input wire spike733,    input wire spike734,    input wire spike735,    input wire spike736,    input wire spike737,    input wire spike738,    input wire spike739,    input wire spike740,    input wire spike741,    input wire spike742,    input wire spike743,    input wire spike744,    input wire spike745,    input wire spike746,    input wire spike747,    input wire spike748,    input wire spike749,    input wire spike750,    input wire spike751,    input wire spike752,    input wire spike753,    input wire spike754,    input wire spike755,    input wire spike756,    input wire spike757,    input wire spike758,    input wire spike759,    input wire spike760,    input wire spike761,    input wire spike762,    input wire spike763,    input wire spike764,    input wire spike765,    input wire spike766,    input wire spike767,    input wire spike768,    input wire spike769,    input wire spike770,    input wire spike771,    input wire spike772,    input wire spike773,    input wire spike774,    input wire spike775,    input wire spike776,    input wire spike777,    input wire spike778,    input wire spike779,    input wire spike780,    input wire spike781,    input wire spike782,    input wire spike783,    input wire spike784,    input wire spike785,    input wire spike786,    input wire spike787,    input wire spike788,    input wire spike789,    input wire spike790,    input wire spike791,    input wire spike792,    input wire spike793,    input wire spike794,    input wire spike795,    input wire spike796,    input wire spike797,    input wire spike798,    input wire spike799,    input wire spike800,
    input wire spike801,    input wire spike802,    input wire spike803,    input wire spike804,    input wire spike805,    input wire spike806,    input wire spike807,    input wire spike808,    input wire spike809,    input wire spike810,    input wire spike811,    input wire spike812,    input wire spike813,    input wire spike814,    input wire spike815,    input wire spike816,    input wire spike817,    input wire spike818,    input wire spike819,    input wire spike820,    input wire spike821,    input wire spike822,    input wire spike823,    input wire spike824,    input wire spike825,    input wire spike826,    input wire spike827,    input wire spike828,    input wire spike829,    input wire spike830,    input wire spike831,    input wire spike832,    input wire spike833,    input wire spike834,    input wire spike835,    input wire spike836,    input wire spike837,    input wire spike838,    input wire spike839,    input wire spike840,    input wire spike841,    input wire spike842,    input wire spike843,    input wire spike844,    input wire spike845,    input wire spike846,    input wire spike847,    input wire spike848,    input wire spike849,    input wire spike850,    input wire spike851,    input wire spike852,    input wire spike853,    input wire spike854,    input wire spike855,    input wire spike856,    input wire spike857,    input wire spike858,    input wire spike859,    input wire spike860,    input wire spike861,    input wire spike862,    input wire spike863,    input wire spike864,    input wire spike865,    input wire spike866,    input wire spike867,    input wire spike868,    input wire spike869,    input wire spike870,    input wire spike871,    input wire spike872,    input wire spike873,    input wire spike874,    input wire spike875,    input wire spike876,    input wire spike877,    input wire spike878,    input wire spike879,    input wire spike880,    input wire spike881,    input wire spike882,    input wire spike883,    input wire spike884,    input wire spike885,    input wire spike886,    input wire spike887,    input wire spike888,    input wire spike889,    input wire spike890,    input wire spike891,    input wire spike892,    input wire spike893,    input wire spike894,    input wire spike895,    input wire spike896,    input wire spike897,    input wire spike898,    input wire spike899,    input wire spike900,
    input wire spike901,    input wire spike902,    input wire spike903,    input wire spike904,    input wire spike905,    input wire spike906,    input wire spike907,    input wire spike908,    input wire spike909,    input wire spike910,    input wire spike911,    input wire spike912,    input wire spike913,    input wire spike914,    input wire spike915,    input wire spike916,    input wire spike917,    input wire spike918,    input wire spike919,    input wire spike920,    input wire spike921,    input wire spike922,    input wire spike923,    input wire spike924,    input wire spike925,    input wire spike926,    input wire spike927,    input wire spike928,    input wire spike929,    input wire spike930,    input wire spike931,    input wire spike932,    input wire spike933,    input wire spike934,    input wire spike935,    input wire spike936,    input wire spike937,    input wire spike938,    input wire spike939,    input wire spike940,    input wire spike941,    input wire spike942,    input wire spike943,    input wire spike944,    input wire spike945,    input wire spike946,    input wire spike947,    input wire spike948,    input wire spike949,    input wire spike950,    input wire spike951,    input wire spike952,    input wire spike953,    input wire spike954,    input wire spike955,    input wire spike956,    input wire spike957,    input wire spike958,    input wire spike959,    input wire spike960,    input wire spike961,    input wire spike962,    input wire spike963,    input wire spike964,    input wire spike965,    input wire spike966,    input wire spike967,    input wire spike968,    input wire spike969,    input wire spike970,    input wire spike971,    input wire spike972,    input wire spike973,    input wire spike974,    input wire spike975,    input wire spike976,    input wire spike977,    input wire spike978,    input wire spike979,    input wire spike980,    input wire spike981,    input wire spike982,    input wire spike983,    input wire spike984,    input wire spike985,    input wire spike986,    input wire spike987,    input wire spike988,    input wire spike989,    input wire spike990,    input wire spike991,    input wire spike992,    input wire spike993,    input wire spike994,    input wire spike995,    input wire spike996,    input wire spike997,    input wire spike998,    input wire spike999,    input wire spike1000,
    input wire spike1001,    input wire spike1002,    input wire spike1003,    input wire spike1004,    input wire spike1005,    input wire spike1006,    input wire spike1007,    input wire spike1008,    input wire spike1009,    input wire spike1010,    input wire spike1011,    input wire spike1012,    input wire spike1013,    input wire spike1014,    input wire spike1015,    input wire spike1016,    input wire spike1017,    input wire spike1018,    input wire spike1019,    input wire spike1020,    input wire spike1021,    input wire spike1022,    input wire spike1023,
output reg[11:0]     spike_out_source0,
    spike_out_source1,    spike_out_source2,    spike_out_source3,    spike_out_source4,    spike_out_source5,    spike_out_source6,    spike_out_source7,    spike_out_source8,    spike_out_source9,    spike_out_source10,    spike_out_source11,    spike_out_source12,    spike_out_source13,    spike_out_source14,    spike_out_source15,    spike_out_source16,    spike_out_source17,    spike_out_source18,    spike_out_source19,    spike_out_source20,    spike_out_source21,    spike_out_source22,    spike_out_source23,    spike_out_source24,    spike_out_source25,    spike_out_source26,    spike_out_source27,    spike_out_source28,    spike_out_source29,    spike_out_source30,    spike_out_source31,    spike_out_source32,    spike_out_source33,    spike_out_source34,    spike_out_source35,    spike_out_source36,    spike_out_source37,    spike_out_source38,    spike_out_source39,    spike_out_source40,    spike_out_source41,    spike_out_source42,    spike_out_source43,    spike_out_source44,    spike_out_source45,    spike_out_source46,    spike_out_source47,    spike_out_source48,    spike_out_source49,    spike_out_source50,    spike_out_source51,    spike_out_source52,    spike_out_source53,    spike_out_source54,    spike_out_source55,    spike_out_source56,    spike_out_source57,    spike_out_source58,    spike_out_source59,    spike_out_source60,    spike_out_source61,    spike_out_source62,    spike_out_source63,    spike_out_source64,    spike_out_source65,    spike_out_source66,    spike_out_source67,    spike_out_source68,    spike_out_source69,    spike_out_source70,    spike_out_source71,    spike_out_source72,    spike_out_source73,    spike_out_source74,    spike_out_source75,    spike_out_source76,    spike_out_source77,    spike_out_source78,    spike_out_source79,    spike_out_source80,    spike_out_source81,    spike_out_source82,    spike_out_source83,    spike_out_source84,    spike_out_source85,    spike_out_source86,    spike_out_source87,    spike_out_source88,    spike_out_source89,    spike_out_source90,    spike_out_source91,    spike_out_source92,    spike_out_source93,    spike_out_source94,    spike_out_source95,    spike_out_source96,    spike_out_source97,    spike_out_source98,    spike_out_source99,    spike_out_source100,
    spike_out_source101,    spike_out_source102,    spike_out_source103,    spike_out_source104,    spike_out_source105,    spike_out_source106,    spike_out_source107,    spike_out_source108,    spike_out_source109,    spike_out_source110,    spike_out_source111,    spike_out_source112,    spike_out_source113,    spike_out_source114,    spike_out_source115,    spike_out_source116,    spike_out_source117,    spike_out_source118,    spike_out_source119,    spike_out_source120,    spike_out_source121,    spike_out_source122,    spike_out_source123,    spike_out_source124,    spike_out_source125,    spike_out_source126,    spike_out_source127,    spike_out_source128,    spike_out_source129,    spike_out_source130,    spike_out_source131,    spike_out_source132,    spike_out_source133,    spike_out_source134,    spike_out_source135,    spike_out_source136,    spike_out_source137,    spike_out_source138,    spike_out_source139,    spike_out_source140,    spike_out_source141,    spike_out_source142,    spike_out_source143,    spike_out_source144,    spike_out_source145,    spike_out_source146,    spike_out_source147,    spike_out_source148,    spike_out_source149,    spike_out_source150,    spike_out_source151,    spike_out_source152,    spike_out_source153,    spike_out_source154,    spike_out_source155,    spike_out_source156,    spike_out_source157,    spike_out_source158,    spike_out_source159,    spike_out_source160,    spike_out_source161,    spike_out_source162,    spike_out_source163,    spike_out_source164,    spike_out_source165,    spike_out_source166,    spike_out_source167,    spike_out_source168,    spike_out_source169,    spike_out_source170,    spike_out_source171,    spike_out_source172,    spike_out_source173,    spike_out_source174,    spike_out_source175,    spike_out_source176,    spike_out_source177,    spike_out_source178,    spike_out_source179,    spike_out_source180,    spike_out_source181,    spike_out_source182,    spike_out_source183,    spike_out_source184,    spike_out_source185,    spike_out_source186,    spike_out_source187,    spike_out_source188,    spike_out_source189,    spike_out_source190,    spike_out_source191,    spike_out_source192,    spike_out_source193,    spike_out_source194,    spike_out_source195,    spike_out_source196,    spike_out_source197,    spike_out_source198,    spike_out_source199,    spike_out_source200,
    spike_out_source201,    spike_out_source202,    spike_out_source203,    spike_out_source204,    spike_out_source205,    spike_out_source206,    spike_out_source207,    spike_out_source208,    spike_out_source209,    spike_out_source210,    spike_out_source211,    spike_out_source212,    spike_out_source213,    spike_out_source214,    spike_out_source215,    spike_out_source216,    spike_out_source217,    spike_out_source218,    spike_out_source219,    spike_out_source220,    spike_out_source221,    spike_out_source222,    spike_out_source223,    spike_out_source224,    spike_out_source225,    spike_out_source226,    spike_out_source227,    spike_out_source228,    spike_out_source229,    spike_out_source230,    spike_out_source231,    spike_out_source232,    spike_out_source233,    spike_out_source234,    spike_out_source235,    spike_out_source236,    spike_out_source237,    spike_out_source238,    spike_out_source239,    spike_out_source240,    spike_out_source241,    spike_out_source242,    spike_out_source243,    spike_out_source244,    spike_out_source245,    spike_out_source246,    spike_out_source247,    spike_out_source248,    spike_out_source249,    spike_out_source250,    spike_out_source251,    spike_out_source252,    spike_out_source253,    spike_out_source254,    spike_out_source255,    spike_out_source256,    spike_out_source257,    spike_out_source258,    spike_out_source259,    spike_out_source260,    spike_out_source261,    spike_out_source262,    spike_out_source263,    spike_out_source264,    spike_out_source265,    spike_out_source266,    spike_out_source267,    spike_out_source268,    spike_out_source269,    spike_out_source270,    spike_out_source271,    spike_out_source272,    spike_out_source273,    spike_out_source274,    spike_out_source275,    spike_out_source276,    spike_out_source277,    spike_out_source278,    spike_out_source279,    spike_out_source280,    spike_out_source281,    spike_out_source282,    spike_out_source283,    spike_out_source284,    spike_out_source285,    spike_out_source286,    spike_out_source287,    spike_out_source288,    spike_out_source289,    spike_out_source290,    spike_out_source291,    spike_out_source292,    spike_out_source293,    spike_out_source294,    spike_out_source295,    spike_out_source296,    spike_out_source297,    spike_out_source298,    spike_out_source299,    spike_out_source300,
    spike_out_source301,    spike_out_source302,    spike_out_source303,    spike_out_source304,    spike_out_source305,    spike_out_source306,    spike_out_source307,    spike_out_source308,    spike_out_source309,    spike_out_source310,    spike_out_source311,    spike_out_source312,    spike_out_source313,    spike_out_source314,    spike_out_source315,    spike_out_source316,    spike_out_source317,    spike_out_source318,    spike_out_source319,    spike_out_source320,    spike_out_source321,    spike_out_source322,    spike_out_source323,    spike_out_source324,    spike_out_source325,    spike_out_source326,    spike_out_source327,    spike_out_source328,    spike_out_source329,    spike_out_source330,    spike_out_source331,    spike_out_source332,    spike_out_source333,    spike_out_source334,    spike_out_source335,    spike_out_source336,    spike_out_source337,    spike_out_source338,    spike_out_source339,    spike_out_source340,    spike_out_source341,    spike_out_source342,    spike_out_source343,    spike_out_source344,    spike_out_source345,    spike_out_source346,    spike_out_source347,    spike_out_source348,    spike_out_source349,    spike_out_source350,    spike_out_source351,    spike_out_source352,    spike_out_source353,    spike_out_source354,    spike_out_source355,    spike_out_source356,    spike_out_source357,    spike_out_source358,    spike_out_source359,    spike_out_source360,    spike_out_source361,    spike_out_source362,    spike_out_source363,    spike_out_source364,    spike_out_source365,    spike_out_source366,    spike_out_source367,    spike_out_source368,    spike_out_source369,    spike_out_source370,    spike_out_source371,    spike_out_source372,    spike_out_source373,    spike_out_source374,    spike_out_source375,    spike_out_source376,    spike_out_source377,    spike_out_source378,    spike_out_source379,    spike_out_source380,    spike_out_source381,    spike_out_source382,    spike_out_source383,    spike_out_source384,    spike_out_source385,    spike_out_source386,    spike_out_source387,    spike_out_source388,    spike_out_source389,    spike_out_source390,    spike_out_source391,    spike_out_source392,    spike_out_source393,    spike_out_source394,    spike_out_source395,    spike_out_source396,    spike_out_source397,    spike_out_source398,    spike_out_source399,    spike_out_source400,
    spike_out_source401,    spike_out_source402,    spike_out_source403,    spike_out_source404,    spike_out_source405,    spike_out_source406,    spike_out_source407,    spike_out_source408,    spike_out_source409,    spike_out_source410,    spike_out_source411,    spike_out_source412,    spike_out_source413,    spike_out_source414,    spike_out_source415,    spike_out_source416,    spike_out_source417,    spike_out_source418,    spike_out_source419,    spike_out_source420,    spike_out_source421,    spike_out_source422,    spike_out_source423,    spike_out_source424,    spike_out_source425,    spike_out_source426,    spike_out_source427,    spike_out_source428,    spike_out_source429,    spike_out_source430,    spike_out_source431,    spike_out_source432,    spike_out_source433,    spike_out_source434,    spike_out_source435,    spike_out_source436,    spike_out_source437,    spike_out_source438,    spike_out_source439,    spike_out_source440,    spike_out_source441,    spike_out_source442,    spike_out_source443,    spike_out_source444,    spike_out_source445,    spike_out_source446,    spike_out_source447,    spike_out_source448,    spike_out_source449,    spike_out_source450,    spike_out_source451,    spike_out_source452,    spike_out_source453,    spike_out_source454,    spike_out_source455,    spike_out_source456,    spike_out_source457,    spike_out_source458,    spike_out_source459,    spike_out_source460,    spike_out_source461,    spike_out_source462,    spike_out_source463,    spike_out_source464,    spike_out_source465,    spike_out_source466,    spike_out_source467,    spike_out_source468,    spike_out_source469,    spike_out_source470,    spike_out_source471,    spike_out_source472,    spike_out_source473,    spike_out_source474,    spike_out_source475,    spike_out_source476,    spike_out_source477,    spike_out_source478,    spike_out_source479,    spike_out_source480,    spike_out_source481,    spike_out_source482,    spike_out_source483,    spike_out_source484,    spike_out_source485,    spike_out_source486,    spike_out_source487,    spike_out_source488,    spike_out_source489,    spike_out_source490,    spike_out_source491,    spike_out_source492,    spike_out_source493,    spike_out_source494,    spike_out_source495,    spike_out_source496,    spike_out_source497,    spike_out_source498,    spike_out_source499,    spike_out_source500,
    spike_out_source501,    spike_out_source502,    spike_out_source503,    spike_out_source504,    spike_out_source505,    spike_out_source506,    spike_out_source507,    spike_out_source508,    spike_out_source509,    spike_out_source510,    spike_out_source511,    spike_out_source512,    spike_out_source513,    spike_out_source514,    spike_out_source515,    spike_out_source516,    spike_out_source517,    spike_out_source518,    spike_out_source519,    spike_out_source520,    spike_out_source521,    spike_out_source522,    spike_out_source523,    spike_out_source524,    spike_out_source525,    spike_out_source526,    spike_out_source527,    spike_out_source528,    spike_out_source529,    spike_out_source530,    spike_out_source531,    spike_out_source532,    spike_out_source533,    spike_out_source534,    spike_out_source535,    spike_out_source536,    spike_out_source537,    spike_out_source538,    spike_out_source539,    spike_out_source540,    spike_out_source541,    spike_out_source542,    spike_out_source543,    spike_out_source544,    spike_out_source545,    spike_out_source546,    spike_out_source547,    spike_out_source548,    spike_out_source549,    spike_out_source550,    spike_out_source551,    spike_out_source552,    spike_out_source553,    spike_out_source554,    spike_out_source555,    spike_out_source556,    spike_out_source557,    spike_out_source558,    spike_out_source559,    spike_out_source560,    spike_out_source561,    spike_out_source562,    spike_out_source563,    spike_out_source564,    spike_out_source565,    spike_out_source566,    spike_out_source567,    spike_out_source568,    spike_out_source569,    spike_out_source570,    spike_out_source571,    spike_out_source572,    spike_out_source573,    spike_out_source574,    spike_out_source575,    spike_out_source576,    spike_out_source577,    spike_out_source578,    spike_out_source579,    spike_out_source580,    spike_out_source581,    spike_out_source582,    spike_out_source583,    spike_out_source584,    spike_out_source585,    spike_out_source586,    spike_out_source587,    spike_out_source588,    spike_out_source589,    spike_out_source590,    spike_out_source591,    spike_out_source592,    spike_out_source593,    spike_out_source594,    spike_out_source595,    spike_out_source596,    spike_out_source597,    spike_out_source598,    spike_out_source599,    spike_out_source600,
    spike_out_source601,    spike_out_source602,    spike_out_source603,    spike_out_source604,    spike_out_source605,    spike_out_source606,    spike_out_source607,    spike_out_source608,    spike_out_source609,    spike_out_source610,    spike_out_source611,    spike_out_source612,    spike_out_source613,    spike_out_source614,    spike_out_source615,    spike_out_source616,    spike_out_source617,    spike_out_source618,    spike_out_source619,    spike_out_source620,    spike_out_source621,    spike_out_source622,    spike_out_source623,    spike_out_source624,    spike_out_source625,    spike_out_source626,    spike_out_source627,    spike_out_source628,    spike_out_source629,    spike_out_source630,    spike_out_source631,    spike_out_source632,    spike_out_source633,    spike_out_source634,    spike_out_source635,    spike_out_source636,    spike_out_source637,    spike_out_source638,    spike_out_source639,    spike_out_source640,    spike_out_source641,    spike_out_source642,    spike_out_source643,    spike_out_source644,    spike_out_source645,    spike_out_source646,    spike_out_source647,    spike_out_source648,    spike_out_source649,    spike_out_source650,    spike_out_source651,    spike_out_source652,    spike_out_source653,    spike_out_source654,    spike_out_source655,    spike_out_source656,    spike_out_source657,    spike_out_source658,    spike_out_source659,    spike_out_source660,    spike_out_source661,    spike_out_source662,    spike_out_source663,    spike_out_source664,    spike_out_source665,    spike_out_source666,    spike_out_source667,    spike_out_source668,    spike_out_source669,    spike_out_source670,    spike_out_source671,    spike_out_source672,    spike_out_source673,    spike_out_source674,    spike_out_source675,    spike_out_source676,    spike_out_source677,    spike_out_source678,    spike_out_source679,    spike_out_source680,    spike_out_source681,    spike_out_source682,    spike_out_source683,    spike_out_source684,    spike_out_source685,    spike_out_source686,    spike_out_source687,    spike_out_source688,    spike_out_source689,    spike_out_source690,    spike_out_source691,    spike_out_source692,    spike_out_source693,    spike_out_source694,    spike_out_source695,    spike_out_source696,    spike_out_source697,    spike_out_source698,    spike_out_source699,    spike_out_source700,
    spike_out_source701,    spike_out_source702,    spike_out_source703,    spike_out_source704,    spike_out_source705,    spike_out_source706,    spike_out_source707,    spike_out_source708,    spike_out_source709,    spike_out_source710,    spike_out_source711,    spike_out_source712,    spike_out_source713,    spike_out_source714,    spike_out_source715,    spike_out_source716,    spike_out_source717,    spike_out_source718,    spike_out_source719,    spike_out_source720,    spike_out_source721,    spike_out_source722,    spike_out_source723,    spike_out_source724,    spike_out_source725,    spike_out_source726,    spike_out_source727,    spike_out_source728,    spike_out_source729,    spike_out_source730,    spike_out_source731,    spike_out_source732,    spike_out_source733,    spike_out_source734,    spike_out_source735,    spike_out_source736,    spike_out_source737,    spike_out_source738,    spike_out_source739,    spike_out_source740,    spike_out_source741,    spike_out_source742,    spike_out_source743,    spike_out_source744,    spike_out_source745,    spike_out_source746,    spike_out_source747,    spike_out_source748,    spike_out_source749,    spike_out_source750,    spike_out_source751,    spike_out_source752,    spike_out_source753,    spike_out_source754,    spike_out_source755,    spike_out_source756,    spike_out_source757,    spike_out_source758,    spike_out_source759,    spike_out_source760,    spike_out_source761,    spike_out_source762,    spike_out_source763,    spike_out_source764,    spike_out_source765,    spike_out_source766,    spike_out_source767,    spike_out_source768,    spike_out_source769,    spike_out_source770,    spike_out_source771,    spike_out_source772,    spike_out_source773,    spike_out_source774,    spike_out_source775,    spike_out_source776,    spike_out_source777,    spike_out_source778,    spike_out_source779,    spike_out_source780,    spike_out_source781,    spike_out_source782,    spike_out_source783,    spike_out_source784,    spike_out_source785,    spike_out_source786,    spike_out_source787,    spike_out_source788,    spike_out_source789,    spike_out_source790,    spike_out_source791,    spike_out_source792,    spike_out_source793,    spike_out_source794,    spike_out_source795,    spike_out_source796,    spike_out_source797,    spike_out_source798,    spike_out_source799,    spike_out_source800,
    spike_out_source801,    spike_out_source802,    spike_out_source803,    spike_out_source804,    spike_out_source805,    spike_out_source806,    spike_out_source807,    spike_out_source808,    spike_out_source809,    spike_out_source810,    spike_out_source811,    spike_out_source812,    spike_out_source813,    spike_out_source814,    spike_out_source815,    spike_out_source816,    spike_out_source817,    spike_out_source818,    spike_out_source819,    spike_out_source820,    spike_out_source821,    spike_out_source822,    spike_out_source823,    spike_out_source824,    spike_out_source825,    spike_out_source826,    spike_out_source827,    spike_out_source828,    spike_out_source829,    spike_out_source830,    spike_out_source831,    spike_out_source832,    spike_out_source833,    spike_out_source834,    spike_out_source835,    spike_out_source836,    spike_out_source837,    spike_out_source838,    spike_out_source839,    spike_out_source840,    spike_out_source841,    spike_out_source842,    spike_out_source843,    spike_out_source844,    spike_out_source845,    spike_out_source846,    spike_out_source847,    spike_out_source848,    spike_out_source849,    spike_out_source850,    spike_out_source851,    spike_out_source852,    spike_out_source853,    spike_out_source854,    spike_out_source855,    spike_out_source856,    spike_out_source857,    spike_out_source858,    spike_out_source859,    spike_out_source860,    spike_out_source861,    spike_out_source862,    spike_out_source863,    spike_out_source864,    spike_out_source865,    spike_out_source866,    spike_out_source867,    spike_out_source868,    spike_out_source869,    spike_out_source870,    spike_out_source871,    spike_out_source872,    spike_out_source873,    spike_out_source874,    spike_out_source875,    spike_out_source876,    spike_out_source877,    spike_out_source878,    spike_out_source879,    spike_out_source880,    spike_out_source881,    spike_out_source882,    spike_out_source883,    spike_out_source884,    spike_out_source885,    spike_out_source886,    spike_out_source887,    spike_out_source888,    spike_out_source889,    spike_out_source890,    spike_out_source891,    spike_out_source892,    spike_out_source893,    spike_out_source894,    spike_out_source895,    spike_out_source896,    spike_out_source897,    spike_out_source898,    spike_out_source899,    spike_out_source900,
    spike_out_source901,    spike_out_source902,    spike_out_source903,    spike_out_source904,    spike_out_source905,    spike_out_source906,    spike_out_source907,    spike_out_source908,    spike_out_source909,    spike_out_source910,    spike_out_source911,    spike_out_source912,    spike_out_source913,    spike_out_source914,    spike_out_source915,    spike_out_source916,    spike_out_source917,    spike_out_source918,    spike_out_source919,    spike_out_source920,    spike_out_source921,    spike_out_source922,    spike_out_source923,    spike_out_source924,    spike_out_source925,    spike_out_source926,    spike_out_source927,    spike_out_source928,    spike_out_source929,    spike_out_source930,    spike_out_source931,    spike_out_source932,    spike_out_source933,    spike_out_source934,    spike_out_source935,    spike_out_source936,    spike_out_source937,    spike_out_source938,    spike_out_source939,    spike_out_source940,    spike_out_source941,    spike_out_source942,    spike_out_source943,    spike_out_source944,    spike_out_source945,    spike_out_source946,    spike_out_source947,    spike_out_source948,    spike_out_source949,    spike_out_source950,    spike_out_source951,    spike_out_source952,    spike_out_source953,    spike_out_source954,    spike_out_source955,    spike_out_source956,    spike_out_source957,    spike_out_source958,    spike_out_source959,    spike_out_source960,    spike_out_source961,    spike_out_source962,    spike_out_source963,    spike_out_source964,    spike_out_source965,    spike_out_source966,    spike_out_source967,    spike_out_source968,    spike_out_source969,    spike_out_source970,    spike_out_source971,    spike_out_source972,    spike_out_source973,    spike_out_source974,    spike_out_source975,    spike_out_source976,    spike_out_source977,    spike_out_source978,    spike_out_source979,    spike_out_source980,    spike_out_source981,    spike_out_source982,    spike_out_source983,    spike_out_source984,    spike_out_source985,    spike_out_source986,    spike_out_source987,    spike_out_source988,    spike_out_source989,    spike_out_source990,    spike_out_source991,    spike_out_source992,    spike_out_source993,    spike_out_source994,    spike_out_source995,    spike_out_source996,    spike_out_source997,    spike_out_source998,    spike_out_source999,    spike_out_source1000,
    spike_out_source1001,    spike_out_source1002,    spike_out_source1003,    spike_out_source1004,    spike_out_source1005,    spike_out_source1006,    spike_out_source1007,    spike_out_source1008,    spike_out_source1009,    spike_out_source1010,    spike_out_source1011,    spike_out_source1012,    spike_out_source1013,    spike_out_source1014,    spike_out_source1015,    spike_out_source1016,    spike_out_source1017,    spike_out_source1018,    spike_out_source1019,    spike_out_source1020,    spike_out_source1021,    spike_out_source1022,    spike_out_source1023,
    output wire output
);

    parameter number_of_neurons= 1024;
    reg spike_register[0:number_of_neurons-1];
    always @(clear, lock1, spike0, spike1, spike2, spike3, spike4, spike5, spike6, spike7, spike8, spike9, spike10, spike11, spike12, spike13, spike14, spike15, spike16, spike17, spike18, spike19, spike20, spike21, spike22, spike23, spike24, spike25, spike26, spike27, spike28, spike29, spike30, spike31, spike32, spike33, spike34, spike35, spike36, spike37, spike38, spike39, spike40, spike41, spike42, spike43, spike44, spike45, spike46, spike47, spike48, spike49) begin
        spike_register[0] = spike0;

        spike_register[1] = spike1;        spike_register[2] = spike2;        spike_register[3] = spike3;        spike_register[4] = spike4;        spike_register[5] = spike5;        spike_register[6] = spike6;        spike_register[7] = spike7;        spike_register[8] = spike8;        spike_register[9] = spike9;        spike_register[10] = spike10;        spike_register[11] = spike11;        spike_register[12] = spike12;        spike_register[13] = spike13;        spike_register[14] = spike14;        spike_register[15] = spike15;        spike_register[16] = spike16;        spike_register[17] = spike17;        spike_register[18] = spike18;        spike_register[19] = spike19;        spike_register[20] = spike20;        spike_register[21] = spike21;        spike_register[22] = spike22;        spike_register[23] = spike23;        spike_register[24] = spike24;        spike_register[25] = spike25;        spike_register[26] = spike26;        spike_register[27] = spike27;        spike_register[28] = spike28;        spike_register[29] = spike29;        spike_register[30] = spike30;        spike_register[31] = spike31;        spike_register[32] = spike32;        spike_register[33] = spike33;        spike_register[34] = spike34;        spike_register[35] = spike35;        spike_register[36] = spike36;        spike_register[37] = spike37;        spike_register[38] = spike38;        spike_register[39] = spike39;        spike_register[40] = spike40;        spike_register[41] = spike41;        spike_register[42] = spike42;        spike_register[43] = spike43;        spike_register[44] = spike44;        spike_register[45] = spike45;        spike_register[46] = spike46;        spike_register[47] = spike47;        spike_register[48] = spike48;        spike_register[49] = spike49;
        #0.5
        if(clear == 1'b0) begin
            for(i1 = 0; i1 <=49; i1= i1+1) begin
                if(spike_register[i1] == 1 && lock1 == 0) begin
                    lock1 = 1;
                    for(j1 = connection_pointer[i1]; j1 < connection_pointer[i1+1]; j1= j1+1) begin
                        packet1 = #0.1 {neuron_addresses[i1], downstream_connections[j1]};
                    end
                    spike_register[i1] = 0;
                    lock1 = 0;
                end
            end
        end

    end
    always @(clear, lock2, spike50, spike51, spike52, spike53, spike54, spike55, spike56, spike57, spike58, spike59, spike60, spike61, spike62, spike63, spike64, spike65, spike66, spike67, spike68, spike69, spike70, spike71, spike72, spike73, spike74, spike75, spike76, spike77, spike78, spike79, spike80, spike81, spike82, spike83, spike84, spike85, spike86, spike87, spike88, spike89, spike90, spike91, spike92, spike93, spike94, spike95, spike96, spike97, spike98, spike99) begin
        spike_register[50] = spike50;        spike_register[51] = spike51;        spike_register[52] = spike52;        spike_register[53] = spike53;        spike_register[54] = spike54;        spike_register[55] = spike55;        spike_register[56] = spike56;        spike_register[57] = spike57;        spike_register[58] = spike58;        spike_register[59] = spike59;        spike_register[60] = spike60;        spike_register[61] = spike61;        spike_register[62] = spike62;        spike_register[63] = spike63;        spike_register[64] = spike64;        spike_register[65] = spike65;        spike_register[66] = spike66;        spike_register[67] = spike67;        spike_register[68] = spike68;        spike_register[69] = spike69;        spike_register[70] = spike70;        spike_register[71] = spike71;        spike_register[72] = spike72;        spike_register[73] = spike73;        spike_register[74] = spike74;        spike_register[75] = spike75;        spike_register[76] = spike76;        spike_register[77] = spike77;        spike_register[78] = spike78;        spike_register[79] = spike79;        spike_register[80] = spike80;        spike_register[81] = spike81;        spike_register[82] = spike82;        spike_register[83] = spike83;        spike_register[84] = spike84;        spike_register[85] = spike85;        spike_register[86] = spike86;        spike_register[87] = spike87;        spike_register[88] = spike88;        spike_register[89] = spike89;        spike_register[90] = spike90;        spike_register[91] = spike91;        spike_register[92] = spike92;        spike_register[93] = spike93;        spike_register[94] = spike94;        spike_register[95] = spike95;        spike_register[96] = spike96;        spike_register[97] = spike97;        spike_register[98] = spike98;        spike_register[99] = spike99;
        #0.5
        if(clear == 1'b0) begin
            for(i2 = 50; i2 <=99; i2= i2+1) begin
                if(spike_register[i2] == 1 && lock2 == 0) begin
                    lock2 = 1;
                    for(j2 = connection_pointer[i2]; j2 < connection_pointer[i2+1]; j2= j2+1) begin
                        packet2 = #0.1 {neuron_addresses[i2], downstream_connections[j2]};
                    end
                    spike_register[i2] = 0;
                    lock2 = 0;
                end
            end
        end

    end
    always @(clear, lock3, spike100, spike101, spike102, spike103, spike104, spike105, spike106, spike107, spike108, spike109, spike110, spike111, spike112, spike113, spike114, spike115, spike116, spike117, spike118, spike119, spike120, spike121, spike122, spike123, spike124, spike125, spike126, spike127, spike128, spike129, spike130, spike131, spike132, spike133, spike134, spike135, spike136, spike137, spike138, spike139, spike140, spike141, spike142, spike143, spike144, spike145, spike146, spike147, spike148, spike149) begin
        spike_register[100] = spike100;

        spike_register[101] = spike101;        spike_register[102] = spike102;        spike_register[103] = spike103;        spike_register[104] = spike104;        spike_register[105] = spike105;        spike_register[106] = spike106;        spike_register[107] = spike107;        spike_register[108] = spike108;        spike_register[109] = spike109;        spike_register[110] = spike110;        spike_register[111] = spike111;        spike_register[112] = spike112;        spike_register[113] = spike113;        spike_register[114] = spike114;        spike_register[115] = spike115;        spike_register[116] = spike116;        spike_register[117] = spike117;        spike_register[118] = spike118;        spike_register[119] = spike119;        spike_register[120] = spike120;        spike_register[121] = spike121;        spike_register[122] = spike122;        spike_register[123] = spike123;        spike_register[124] = spike124;        spike_register[125] = spike125;        spike_register[126] = spike126;        spike_register[127] = spike127;        spike_register[128] = spike128;        spike_register[129] = spike129;        spike_register[130] = spike130;        spike_register[131] = spike131;        spike_register[132] = spike132;        spike_register[133] = spike133;        spike_register[134] = spike134;        spike_register[135] = spike135;        spike_register[136] = spike136;        spike_register[137] = spike137;        spike_register[138] = spike138;        spike_register[139] = spike139;        spike_register[140] = spike140;        spike_register[141] = spike141;        spike_register[142] = spike142;        spike_register[143] = spike143;        spike_register[144] = spike144;        spike_register[145] = spike145;        spike_register[146] = spike146;        spike_register[147] = spike147;        spike_register[148] = spike148;        spike_register[149] = spike149;
        #0.5
        if(clear == 1'b0) begin
            for(i3 = 100; i3 <=149; i3= i3+1) begin
                if(spike_register[i3] == 1 && lock3 == 0) begin
                    lock3 = 1;
                    for(j3 = connection_pointer[i3]; j3 < connection_pointer[i3+1]; j3= j3+1) begin
                        packet3 = #0.1 {neuron_addresses[i3], downstream_connections[j3]};
                    end
                    spike_register[i3] = 0;
                    lock3 = 0;
                end
            end
        end

    end
    always @(clear, lock4, spike150, spike151, spike152, spike153, spike154, spike155, spike156, spike157, spike158, spike159, spike160, spike161, spike162, spike163, spike164, spike165, spike166, spike167, spike168, spike169, spike170, spike171, spike172, spike173, spike174, spike175, spike176, spike177, spike178, spike179, spike180, spike181, spike182, spike183, spike184, spike185, spike186, spike187, spike188, spike189, spike190, spike191, spike192, spike193, spike194, spike195, spike196, spike197, spike198, spike199) begin
        spike_register[150] = spike150;        spike_register[151] = spike151;        spike_register[152] = spike152;        spike_register[153] = spike153;        spike_register[154] = spike154;        spike_register[155] = spike155;        spike_register[156] = spike156;        spike_register[157] = spike157;        spike_register[158] = spike158;        spike_register[159] = spike159;        spike_register[160] = spike160;        spike_register[161] = spike161;        spike_register[162] = spike162;        spike_register[163] = spike163;        spike_register[164] = spike164;        spike_register[165] = spike165;        spike_register[166] = spike166;        spike_register[167] = spike167;        spike_register[168] = spike168;        spike_register[169] = spike169;        spike_register[170] = spike170;        spike_register[171] = spike171;        spike_register[172] = spike172;        spike_register[173] = spike173;        spike_register[174] = spike174;        spike_register[175] = spike175;        spike_register[176] = spike176;        spike_register[177] = spike177;        spike_register[178] = spike178;        spike_register[179] = spike179;        spike_register[180] = spike180;        spike_register[181] = spike181;        spike_register[182] = spike182;        spike_register[183] = spike183;        spike_register[184] = spike184;        spike_register[185] = spike185;        spike_register[186] = spike186;        spike_register[187] = spike187;        spike_register[188] = spike188;        spike_register[189] = spike189;        spike_register[190] = spike190;        spike_register[191] = spike191;        spike_register[192] = spike192;        spike_register[193] = spike193;        spike_register[194] = spike194;        spike_register[195] = spike195;        spike_register[196] = spike196;        spike_register[197] = spike197;        spike_register[198] = spike198;        spike_register[199] = spike199;
        #0.5
        if(clear == 1'b0) begin
            for(i4 = 150; i4 <=199; i4= i4+1) begin
                if(spike_register[i4] == 1 && lock4 == 0) begin
                    lock4 = 1;
                    for(j4 = connection_pointer[i4]; j4 < connection_pointer[i4+1]; j4= j4+1) begin
                        packet4 = #0.1 {neuron_addresses[i4], downstream_connections[j4]};
                    end
                    spike_register[i4] = 0;
                    lock4 = 0;
                end
            end
        end

    end
    always @(clear, lock5, spike200, spike201, spike202, spike203, spike204, spike205, spike206, spike207, spike208, spike209, spike210, spike211, spike212, spike213, spike214, spike215, spike216, spike217, spike218, spike219, spike220, spike221, spike222, spike223, spike224, spike225, spike226, spike227, spike228, spike229, spike230, spike231, spike232, spike233, spike234, spike235, spike236, spike237, spike238, spike239, spike240, spike241, spike242, spike243, spike244, spike245, spike246, spike247, spike248, spike249) begin
        spike_register[200] = spike200;

        spike_register[201] = spike201;        spike_register[202] = spike202;        spike_register[203] = spike203;        spike_register[204] = spike204;        spike_register[205] = spike205;        spike_register[206] = spike206;        spike_register[207] = spike207;        spike_register[208] = spike208;        spike_register[209] = spike209;        spike_register[210] = spike210;        spike_register[211] = spike211;        spike_register[212] = spike212;        spike_register[213] = spike213;        spike_register[214] = spike214;        spike_register[215] = spike215;        spike_register[216] = spike216;        spike_register[217] = spike217;        spike_register[218] = spike218;        spike_register[219] = spike219;        spike_register[220] = spike220;        spike_register[221] = spike221;        spike_register[222] = spike222;        spike_register[223] = spike223;        spike_register[224] = spike224;        spike_register[225] = spike225;        spike_register[226] = spike226;        spike_register[227] = spike227;        spike_register[228] = spike228;        spike_register[229] = spike229;        spike_register[230] = spike230;        spike_register[231] = spike231;        spike_register[232] = spike232;        spike_register[233] = spike233;        spike_register[234] = spike234;        spike_register[235] = spike235;        spike_register[236] = spike236;        spike_register[237] = spike237;        spike_register[238] = spike238;        spike_register[239] = spike239;        spike_register[240] = spike240;        spike_register[241] = spike241;        spike_register[242] = spike242;        spike_register[243] = spike243;        spike_register[244] = spike244;        spike_register[245] = spike245;        spike_register[246] = spike246;        spike_register[247] = spike247;        spike_register[248] = spike248;        spike_register[249] = spike249;
        #0.5
        if(clear == 1'b0) begin
            for(i5 = 200; i5 <=249; i5= i5+1) begin
                if(spike_register[i5] == 1 && lock5 == 0) begin
                    lock5 = 1;
                    for(j5 = connection_pointer[i5]; j5 < connection_pointer[i5+1]; j5= j5+1) begin
                        packet5 = #0.1 {neuron_addresses[i5], downstream_connections[j5]};
                    end
                    spike_register[i5] = 0;
                    lock5 = 0;
                end
            end
        end

    end
    always @(clear, lock6, spike250, spike251, spike252, spike253, spike254, spike255, spike256, spike257, spike258, spike259, spike260, spike261, spike262, spike263, spike264, spike265, spike266, spike267, spike268, spike269, spike270, spike271, spike272, spike273, spike274, spike275, spike276, spike277, spike278, spike279, spike280, spike281, spike282, spike283, spike284, spike285, spike286, spike287, spike288, spike289, spike290, spike291, spike292, spike293, spike294, spike295, spike296, spike297, spike298, spike299) begin
        spike_register[250] = spike250;        spike_register[251] = spike251;        spike_register[252] = spike252;        spike_register[253] = spike253;        spike_register[254] = spike254;        spike_register[255] = spike255;        spike_register[256] = spike256;        spike_register[257] = spike257;        spike_register[258] = spike258;        spike_register[259] = spike259;        spike_register[260] = spike260;        spike_register[261] = spike261;        spike_register[262] = spike262;        spike_register[263] = spike263;        spike_register[264] = spike264;        spike_register[265] = spike265;        spike_register[266] = spike266;        spike_register[267] = spike267;        spike_register[268] = spike268;        spike_register[269] = spike269;        spike_register[270] = spike270;        spike_register[271] = spike271;        spike_register[272] = spike272;        spike_register[273] = spike273;        spike_register[274] = spike274;        spike_register[275] = spike275;        spike_register[276] = spike276;        spike_register[277] = spike277;        spike_register[278] = spike278;        spike_register[279] = spike279;        spike_register[280] = spike280;        spike_register[281] = spike281;        spike_register[282] = spike282;        spike_register[283] = spike283;        spike_register[284] = spike284;        spike_register[285] = spike285;        spike_register[286] = spike286;        spike_register[287] = spike287;        spike_register[288] = spike288;        spike_register[289] = spike289;        spike_register[290] = spike290;        spike_register[291] = spike291;        spike_register[292] = spike292;        spike_register[293] = spike293;        spike_register[294] = spike294;        spike_register[295] = spike295;        spike_register[296] = spike296;        spike_register[297] = spike297;        spike_register[298] = spike298;        spike_register[299] = spike299;
        #0.5
        if(clear == 1'b0) begin
            for(i6 = 250; i6 <=299; i6= i6+1) begin
                if(spike_register[i6] == 1 && lock6 == 0) begin
                    lock6 = 1;
                    for(j6 = connection_pointer[i6]; j6 < connection_pointer[i6+1]; j6= j6+1) begin
                        packet6 = #0.1 {neuron_addresses[i6], downstream_connections[j6]};
                    end
                    spike_register[i6] = 0;
                    lock6 = 0;
                end
            end
        end

    end
    always @(clear, lock7, spike300, spike301, spike302, spike303, spike304, spike305, spike306, spike307, spike308, spike309, spike310, spike311, spike312, spike313, spike314, spike315, spike316, spike317, spike318, spike319, spike320, spike321, spike322, spike323, spike324, spike325, spike326, spike327, spike328, spike329, spike330, spike331, spike332, spike333, spike334, spike335, spike336, spike337, spike338, spike339, spike340, spike341, spike342, spike343, spike344, spike345, spike346, spike347, spike348, spike349) begin
        spike_register[300] = spike300;

        spike_register[301] = spike301;        spike_register[302] = spike302;        spike_register[303] = spike303;        spike_register[304] = spike304;        spike_register[305] = spike305;        spike_register[306] = spike306;        spike_register[307] = spike307;        spike_register[308] = spike308;        spike_register[309] = spike309;        spike_register[310] = spike310;        spike_register[311] = spike311;        spike_register[312] = spike312;        spike_register[313] = spike313;        spike_register[314] = spike314;        spike_register[315] = spike315;        spike_register[316] = spike316;        spike_register[317] = spike317;        spike_register[318] = spike318;        spike_register[319] = spike319;        spike_register[320] = spike320;        spike_register[321] = spike321;        spike_register[322] = spike322;        spike_register[323] = spike323;        spike_register[324] = spike324;        spike_register[325] = spike325;        spike_register[326] = spike326;        spike_register[327] = spike327;        spike_register[328] = spike328;        spike_register[329] = spike329;        spike_register[330] = spike330;        spike_register[331] = spike331;        spike_register[332] = spike332;        spike_register[333] = spike333;        spike_register[334] = spike334;        spike_register[335] = spike335;        spike_register[336] = spike336;        spike_register[337] = spike337;        spike_register[338] = spike338;        spike_register[339] = spike339;        spike_register[340] = spike340;        spike_register[341] = spike341;        spike_register[342] = spike342;        spike_register[343] = spike343;        spike_register[344] = spike344;        spike_register[345] = spike345;        spike_register[346] = spike346;        spike_register[347] = spike347;        spike_register[348] = spike348;        spike_register[349] = spike349;
        #0.5
        if(clear == 1'b0) begin
            for(i7 = 300; i7 <=349; i7= i7+1) begin
                if(spike_register[i7] == 1 && lock7 == 0) begin
                    lock7 = 1;
                    for(j7 = connection_pointer[i7]; j7 < connection_pointer[i7+1]; j7= j7+1) begin
                        packet7 = #0.1 {neuron_addresses[i7], downstream_connections[j7]};
                    end
                    spike_register[i7] = 0;
                    lock7 = 0;
                end
            end
        end

    end
    always @(clear, lock8, spike350, spike351, spike352, spike353, spike354, spike355, spike356, spike357, spike358, spike359, spike360, spike361, spike362, spike363, spike364, spike365, spike366, spike367, spike368, spike369, spike370, spike371, spike372, spike373, spike374, spike375, spike376, spike377, spike378, spike379, spike380, spike381, spike382, spike383, spike384, spike385, spike386, spike387, spike388, spike389, spike390, spike391, spike392, spike393, spike394, spike395, spike396, spike397, spike398, spike399) begin
        spike_register[350] = spike350;        spike_register[351] = spike351;        spike_register[352] = spike352;        spike_register[353] = spike353;        spike_register[354] = spike354;        spike_register[355] = spike355;        spike_register[356] = spike356;        spike_register[357] = spike357;        spike_register[358] = spike358;        spike_register[359] = spike359;        spike_register[360] = spike360;        spike_register[361] = spike361;        spike_register[362] = spike362;        spike_register[363] = spike363;        spike_register[364] = spike364;        spike_register[365] = spike365;        spike_register[366] = spike366;        spike_register[367] = spike367;        spike_register[368] = spike368;        spike_register[369] = spike369;        spike_register[370] = spike370;        spike_register[371] = spike371;        spike_register[372] = spike372;        spike_register[373] = spike373;        spike_register[374] = spike374;        spike_register[375] = spike375;        spike_register[376] = spike376;        spike_register[377] = spike377;        spike_register[378] = spike378;        spike_register[379] = spike379;        spike_register[380] = spike380;        spike_register[381] = spike381;        spike_register[382] = spike382;        spike_register[383] = spike383;        spike_register[384] = spike384;        spike_register[385] = spike385;        spike_register[386] = spike386;        spike_register[387] = spike387;        spike_register[388] = spike388;        spike_register[389] = spike389;        spike_register[390] = spike390;        spike_register[391] = spike391;        spike_register[392] = spike392;        spike_register[393] = spike393;        spike_register[394] = spike394;        spike_register[395] = spike395;        spike_register[396] = spike396;        spike_register[397] = spike397;        spike_register[398] = spike398;        spike_register[399] = spike399;
        #0.5
        if(clear == 1'b0) begin
            for(i8 = 350; i8 <=399; i8= i8+1) begin
                if(spike_register[i8] == 1 && lock8 == 0) begin
                    lock8 = 1;
                    for(j8 = connection_pointer[i8]; j8 < connection_pointer[i8+1]; j8= j8+1) begin
                        packet8 = #0.1 {neuron_addresses[i8], downstream_connections[j8]};
                    end
                    spike_register[i8] = 0;
                    lock8 = 0;
                end
            end
        end

    end
    always @(clear, lock9, spike400, spike401, spike402, spike403, spike404, spike405, spike406, spike407, spike408, spike409, spike410, spike411, spike412, spike413, spike414, spike415, spike416, spike417, spike418, spike419, spike420, spike421, spike422, spike423, spike424, spike425, spike426, spike427, spike428, spike429, spike430, spike431, spike432, spike433, spike434, spike435, spike436, spike437, spike438, spike439, spike440, spike441, spike442, spike443, spike444, spike445, spike446, spike447, spike448, spike449) begin
        spike_register[400] = spike400;

        spike_register[401] = spike401;        spike_register[402] = spike402;        spike_register[403] = spike403;        spike_register[404] = spike404;        spike_register[405] = spike405;        spike_register[406] = spike406;        spike_register[407] = spike407;        spike_register[408] = spike408;        spike_register[409] = spike409;        spike_register[410] = spike410;        spike_register[411] = spike411;        spike_register[412] = spike412;        spike_register[413] = spike413;        spike_register[414] = spike414;        spike_register[415] = spike415;        spike_register[416] = spike416;        spike_register[417] = spike417;        spike_register[418] = spike418;        spike_register[419] = spike419;        spike_register[420] = spike420;        spike_register[421] = spike421;        spike_register[422] = spike422;        spike_register[423] = spike423;        spike_register[424] = spike424;        spike_register[425] = spike425;        spike_register[426] = spike426;        spike_register[427] = spike427;        spike_register[428] = spike428;        spike_register[429] = spike429;        spike_register[430] = spike430;        spike_register[431] = spike431;        spike_register[432] = spike432;        spike_register[433] = spike433;        spike_register[434] = spike434;        spike_register[435] = spike435;        spike_register[436] = spike436;        spike_register[437] = spike437;        spike_register[438] = spike438;        spike_register[439] = spike439;        spike_register[440] = spike440;        spike_register[441] = spike441;        spike_register[442] = spike442;        spike_register[443] = spike443;        spike_register[444] = spike444;        spike_register[445] = spike445;        spike_register[446] = spike446;        spike_register[447] = spike447;        spike_register[448] = spike448;        spike_register[449] = spike449;
        #0.5
        if(clear == 1'b0) begin
            for(i9 = 400; i9 <=449; i9= i9+1) begin
                if(spike_register[i9] == 1 && lock9 == 0) begin
                    lock9 = 1;
                    for(j9 = connection_pointer[i9]; j9 < connection_pointer[i9+1]; j9= j9+1) begin
                        packet9 = #0.1 {neuron_addresses[i9], downstream_connections[j9]};
                    end
                    spike_register[i9] = 0;
                    lock9 = 0;
                end
            end
        end

    end
    always @(clear, lock10, spike450, spike451, spike452, spike453, spike454, spike455, spike456, spike457, spike458, spike459, spike460, spike461, spike462, spike463, spike464, spike465, spike466, spike467, spike468, spike469, spike470, spike471, spike472, spike473, spike474, spike475, spike476, spike477, spike478, spike479, spike480, spike481, spike482, spike483, spike484, spike485, spike486, spike487, spike488, spike489, spike490, spike491, spike492, spike493, spike494, spike495, spike496, spike497, spike498, spike499) begin
        spike_register[450] = spike450;        spike_register[451] = spike451;        spike_register[452] = spike452;        spike_register[453] = spike453;        spike_register[454] = spike454;        spike_register[455] = spike455;        spike_register[456] = spike456;        spike_register[457] = spike457;        spike_register[458] = spike458;        spike_register[459] = spike459;        spike_register[460] = spike460;        spike_register[461] = spike461;        spike_register[462] = spike462;        spike_register[463] = spike463;        spike_register[464] = spike464;        spike_register[465] = spike465;        spike_register[466] = spike466;        spike_register[467] = spike467;        spike_register[468] = spike468;        spike_register[469] = spike469;        spike_register[470] = spike470;        spike_register[471] = spike471;        spike_register[472] = spike472;        spike_register[473] = spike473;        spike_register[474] = spike474;        spike_register[475] = spike475;        spike_register[476] = spike476;        spike_register[477] = spike477;        spike_register[478] = spike478;        spike_register[479] = spike479;        spike_register[480] = spike480;        spike_register[481] = spike481;        spike_register[482] = spike482;        spike_register[483] = spike483;        spike_register[484] = spike484;        spike_register[485] = spike485;        spike_register[486] = spike486;        spike_register[487] = spike487;        spike_register[488] = spike488;        spike_register[489] = spike489;        spike_register[490] = spike490;        spike_register[491] = spike491;        spike_register[492] = spike492;        spike_register[493] = spike493;        spike_register[494] = spike494;        spike_register[495] = spike495;        spike_register[496] = spike496;        spike_register[497] = spike497;        spike_register[498] = spike498;        spike_register[499] = spike499;
        #0.5
        if(clear == 1'b0) begin
            for(i10 = 450; i10 <=499; i10= i10+1) begin
                if(spike_register[i10] == 1 && lock10 == 0) begin
                    lock10 = 1;
                    for(j10 = connection_pointer[i10]; j10 < connection_pointer[i10+1]; j10= j10+1) begin
                        packet10 = #0.1 {neuron_addresses[i10], downstream_connections[j10]};
                    end
                    spike_register[i10] = 0;
                    lock10 = 0;
                end
            end
        end

    end
    always @(clear, lock11, spike500, spike501, spike502, spike503, spike504, spike505, spike506, spike507, spike508, spike509, spike510, spike511, spike512, spike513, spike514, spike515, spike516, spike517, spike518, spike519, spike520, spike521, spike522, spike523, spike524, spike525, spike526, spike527, spike528, spike529, spike530, spike531, spike532, spike533, spike534, spike535, spike536, spike537, spike538, spike539, spike540, spike541, spike542, spike543, spike544, spike545, spike546, spike547, spike548, spike549) begin
        spike_register[500] = spike500;

        spike_register[501] = spike501;        spike_register[502] = spike502;        spike_register[503] = spike503;        spike_register[504] = spike504;        spike_register[505] = spike505;        spike_register[506] = spike506;        spike_register[507] = spike507;        spike_register[508] = spike508;        spike_register[509] = spike509;        spike_register[510] = spike510;        spike_register[511] = spike511;        spike_register[512] = spike512;        spike_register[513] = spike513;        spike_register[514] = spike514;        spike_register[515] = spike515;        spike_register[516] = spike516;        spike_register[517] = spike517;        spike_register[518] = spike518;        spike_register[519] = spike519;        spike_register[520] = spike520;        spike_register[521] = spike521;        spike_register[522] = spike522;        spike_register[523] = spike523;        spike_register[524] = spike524;        spike_register[525] = spike525;        spike_register[526] = spike526;        spike_register[527] = spike527;        spike_register[528] = spike528;        spike_register[529] = spike529;        spike_register[530] = spike530;        spike_register[531] = spike531;        spike_register[532] = spike532;        spike_register[533] = spike533;        spike_register[534] = spike534;        spike_register[535] = spike535;        spike_register[536] = spike536;        spike_register[537] = spike537;        spike_register[538] = spike538;        spike_register[539] = spike539;        spike_register[540] = spike540;        spike_register[541] = spike541;        spike_register[542] = spike542;        spike_register[543] = spike543;        spike_register[544] = spike544;        spike_register[545] = spike545;        spike_register[546] = spike546;        spike_register[547] = spike547;        spike_register[548] = spike548;        spike_register[549] = spike549;
        #0.5
        if(clear == 1'b0) begin
            for(i11 = 500; i11 <=549; i11= i11+1) begin
                if(spike_register[i11] == 1 && lock11 == 0) begin
                    lock11 = 1;
                    for(j11 = connection_pointer[i11]; j11 < connection_pointer[i11+1]; j11= j11+1) begin
                        packet11 = #0.1 {neuron_addresses[i11], downstream_connections[j11]};
                    end
                    spike_register[i11] = 0;
                    lock11 = 0;
                end
            end
        end

    end
    always @(clear, lock12, spike550, spike551, spike552, spike553, spike554, spike555, spike556, spike557, spike558, spike559, spike560, spike561, spike562, spike563, spike564, spike565, spike566, spike567, spike568, spike569, spike570, spike571, spike572, spike573, spike574, spike575, spike576, spike577, spike578, spike579, spike580, spike581, spike582, spike583, spike584, spike585, spike586, spike587, spike588, spike589, spike590, spike591, spike592, spike593, spike594, spike595, spike596, spike597, spike598, spike599) begin
        spike_register[550] = spike550;        spike_register[551] = spike551;        spike_register[552] = spike552;        spike_register[553] = spike553;        spike_register[554] = spike554;        spike_register[555] = spike555;        spike_register[556] = spike556;        spike_register[557] = spike557;        spike_register[558] = spike558;        spike_register[559] = spike559;        spike_register[560] = spike560;        spike_register[561] = spike561;        spike_register[562] = spike562;        spike_register[563] = spike563;        spike_register[564] = spike564;        spike_register[565] = spike565;        spike_register[566] = spike566;        spike_register[567] = spike567;        spike_register[568] = spike568;        spike_register[569] = spike569;        spike_register[570] = spike570;        spike_register[571] = spike571;        spike_register[572] = spike572;        spike_register[573] = spike573;        spike_register[574] = spike574;        spike_register[575] = spike575;        spike_register[576] = spike576;        spike_register[577] = spike577;        spike_register[578] = spike578;        spike_register[579] = spike579;        spike_register[580] = spike580;        spike_register[581] = spike581;        spike_register[582] = spike582;        spike_register[583] = spike583;        spike_register[584] = spike584;        spike_register[585] = spike585;        spike_register[586] = spike586;        spike_register[587] = spike587;        spike_register[588] = spike588;        spike_register[589] = spike589;        spike_register[590] = spike590;        spike_register[591] = spike591;        spike_register[592] = spike592;        spike_register[593] = spike593;        spike_register[594] = spike594;        spike_register[595] = spike595;        spike_register[596] = spike596;        spike_register[597] = spike597;        spike_register[598] = spike598;        spike_register[599] = spike599;
        #0.5
        if(clear == 1'b0) begin
            for(i12 = 550; i12 <=599; i12= i12+1) begin
                if(spike_register[i12] == 1 && lock12 == 0) begin
                    lock12 = 1;
                    for(j12 = connection_pointer[i12]; j12 < connection_pointer[i12+1]; j12= j12+1) begin
                        packet12 = #0.1 {neuron_addresses[i12], downstream_connections[j12]};
                    end
                    spike_register[i12] = 0;
                    lock12 = 0;
                end
            end
        end

    end
    always @(clear, lock13, spike600, spike601, spike602, spike603, spike604, spike605, spike606, spike607, spike608, spike609, spike610, spike611, spike612, spike613, spike614, spike615, spike616, spike617, spike618, spike619, spike620, spike621, spike622, spike623, spike624, spike625, spike626, spike627, spike628, spike629, spike630, spike631, spike632, spike633, spike634, spike635, spike636, spike637, spike638, spike639, spike640, spike641, spike642, spike643, spike644, spike645, spike646, spike647, spike648, spike649) begin
        spike_register[600] = spike600;

        spike_register[601] = spike601;        spike_register[602] = spike602;        spike_register[603] = spike603;        spike_register[604] = spike604;        spike_register[605] = spike605;        spike_register[606] = spike606;        spike_register[607] = spike607;        spike_register[608] = spike608;        spike_register[609] = spike609;        spike_register[610] = spike610;        spike_register[611] = spike611;        spike_register[612] = spike612;        spike_register[613] = spike613;        spike_register[614] = spike614;        spike_register[615] = spike615;        spike_register[616] = spike616;        spike_register[617] = spike617;        spike_register[618] = spike618;        spike_register[619] = spike619;        spike_register[620] = spike620;        spike_register[621] = spike621;        spike_register[622] = spike622;        spike_register[623] = spike623;        spike_register[624] = spike624;        spike_register[625] = spike625;        spike_register[626] = spike626;        spike_register[627] = spike627;        spike_register[628] = spike628;        spike_register[629] = spike629;        spike_register[630] = spike630;        spike_register[631] = spike631;        spike_register[632] = spike632;        spike_register[633] = spike633;        spike_register[634] = spike634;        spike_register[635] = spike635;        spike_register[636] = spike636;        spike_register[637] = spike637;        spike_register[638] = spike638;        spike_register[639] = spike639;        spike_register[640] = spike640;        spike_register[641] = spike641;        spike_register[642] = spike642;        spike_register[643] = spike643;        spike_register[644] = spike644;        spike_register[645] = spike645;        spike_register[646] = spike646;        spike_register[647] = spike647;        spike_register[648] = spike648;        spike_register[649] = spike649;
        #0.5
        if(clear == 1'b0) begin
            for(i13 = 600; i13 <=649; i13= i13+1) begin
                if(spike_register[i13] == 1 && lock13 == 0) begin
                    lock13 = 1;
                    for(j13 = connection_pointer[i13]; j13 < connection_pointer[i13+1]; j13= j13+1) begin
                        packet13 = #0.1 {neuron_addresses[i13], downstream_connections[j13]};
                    end
                    spike_register[i13] = 0;
                    lock13 = 0;
                end
            end
        end

    end
    always @(clear, lock14, spike650, spike651, spike652, spike653, spike654, spike655, spike656, spike657, spike658, spike659, spike660, spike661, spike662, spike663, spike664, spike665, spike666, spike667, spike668, spike669, spike670, spike671, spike672, spike673, spike674, spike675, spike676, spike677, spike678, spike679, spike680, spike681, spike682, spike683, spike684, spike685, spike686, spike687, spike688, spike689, spike690, spike691, spike692, spike693, spike694, spike695, spike696, spike697, spike698, spike699) begin
        spike_register[650] = spike650;        spike_register[651] = spike651;        spike_register[652] = spike652;        spike_register[653] = spike653;        spike_register[654] = spike654;        spike_register[655] = spike655;        spike_register[656] = spike656;        spike_register[657] = spike657;        spike_register[658] = spike658;        spike_register[659] = spike659;        spike_register[660] = spike660;        spike_register[661] = spike661;        spike_register[662] = spike662;        spike_register[663] = spike663;        spike_register[664] = spike664;        spike_register[665] = spike665;        spike_register[666] = spike666;        spike_register[667] = spike667;        spike_register[668] = spike668;        spike_register[669] = spike669;        spike_register[670] = spike670;        spike_register[671] = spike671;        spike_register[672] = spike672;        spike_register[673] = spike673;        spike_register[674] = spike674;        spike_register[675] = spike675;        spike_register[676] = spike676;        spike_register[677] = spike677;        spike_register[678] = spike678;        spike_register[679] = spike679;        spike_register[680] = spike680;        spike_register[681] = spike681;        spike_register[682] = spike682;        spike_register[683] = spike683;        spike_register[684] = spike684;        spike_register[685] = spike685;        spike_register[686] = spike686;        spike_register[687] = spike687;        spike_register[688] = spike688;        spike_register[689] = spike689;        spike_register[690] = spike690;        spike_register[691] = spike691;        spike_register[692] = spike692;        spike_register[693] = spike693;        spike_register[694] = spike694;        spike_register[695] = spike695;        spike_register[696] = spike696;        spike_register[697] = spike697;        spike_register[698] = spike698;        spike_register[699] = spike699;
        #0.5
        if(clear == 1'b0) begin
            for(i14 = 650; i14 <=699; i14= i14+1) begin
                if(spike_register[i14] == 1 && lock14 == 0) begin
                    lock14 = 1;
                    for(j14 = connection_pointer[i14]; j14 < connection_pointer[i14+1]; j14= j14+1) begin
                        packet14 = #0.1 {neuron_addresses[i14], downstream_connections[j14]};
                    end
                    spike_register[i14] = 0;
                    lock14 = 0;
                end
            end
        end

    end
    always @(clear, lock15, spike700, spike701, spike702, spike703, spike704, spike705, spike706, spike707, spike708, spike709, spike710, spike711, spike712, spike713, spike714, spike715, spike716, spike717, spike718, spike719, spike720, spike721, spike722, spike723, spike724, spike725, spike726, spike727, spike728, spike729, spike730, spike731, spike732, spike733, spike734, spike735, spike736, spike737, spike738, spike739, spike740, spike741, spike742, spike743, spike744, spike745, spike746, spike747, spike748, spike749) begin
        spike_register[700] = spike700;

        spike_register[701] = spike701;        spike_register[702] = spike702;        spike_register[703] = spike703;        spike_register[704] = spike704;        spike_register[705] = spike705;        spike_register[706] = spike706;        spike_register[707] = spike707;        spike_register[708] = spike708;        spike_register[709] = spike709;        spike_register[710] = spike710;        spike_register[711] = spike711;        spike_register[712] = spike712;        spike_register[713] = spike713;        spike_register[714] = spike714;        spike_register[715] = spike715;        spike_register[716] = spike716;        spike_register[717] = spike717;        spike_register[718] = spike718;        spike_register[719] = spike719;        spike_register[720] = spike720;        spike_register[721] = spike721;        spike_register[722] = spike722;        spike_register[723] = spike723;        spike_register[724] = spike724;        spike_register[725] = spike725;        spike_register[726] = spike726;        spike_register[727] = spike727;        spike_register[728] = spike728;        spike_register[729] = spike729;        spike_register[730] = spike730;        spike_register[731] = spike731;        spike_register[732] = spike732;        spike_register[733] = spike733;        spike_register[734] = spike734;        spike_register[735] = spike735;        spike_register[736] = spike736;        spike_register[737] = spike737;        spike_register[738] = spike738;        spike_register[739] = spike739;        spike_register[740] = spike740;        spike_register[741] = spike741;        spike_register[742] = spike742;        spike_register[743] = spike743;        spike_register[744] = spike744;        spike_register[745] = spike745;        spike_register[746] = spike746;        spike_register[747] = spike747;        spike_register[748] = spike748;        spike_register[749] = spike749;
        #0.5
        if(clear == 1'b0) begin
            for(i15 = 700; i15 <=749; i15= i15+1) begin
                if(spike_register[i15] == 1 && lock15 == 0) begin
                    lock15 = 1;
                    for(j15 = connection_pointer[i15]; j15 < connection_pointer[i15+1]; j15= j15+1) begin
                        packet15 = #0.1 {neuron_addresses[i15], downstream_connections[j15]};
                    end
                    spike_register[i15] = 0;
                    lock15 = 0;
                end
            end
        end

    end
    always @(clear, lock16, spike750, spike751, spike752, spike753, spike754, spike755, spike756, spike757, spike758, spike759, spike760, spike761, spike762, spike763, spike764, spike765, spike766, spike767, spike768, spike769, spike770, spike771, spike772, spike773, spike774, spike775, spike776, spike777, spike778, spike779, spike780, spike781, spike782, spike783, spike784, spike785, spike786, spike787, spike788, spike789, spike790, spike791, spike792, spike793, spike794, spike795, spike796, spike797, spike798, spike799) begin
        spike_register[750] = spike750;        spike_register[751] = spike751;        spike_register[752] = spike752;        spike_register[753] = spike753;        spike_register[754] = spike754;        spike_register[755] = spike755;        spike_register[756] = spike756;        spike_register[757] = spike757;        spike_register[758] = spike758;        spike_register[759] = spike759;        spike_register[760] = spike760;        spike_register[761] = spike761;        spike_register[762] = spike762;        spike_register[763] = spike763;        spike_register[764] = spike764;        spike_register[765] = spike765;        spike_register[766] = spike766;        spike_register[767] = spike767;        spike_register[768] = spike768;        spike_register[769] = spike769;        spike_register[770] = spike770;        spike_register[771] = spike771;        spike_register[772] = spike772;        spike_register[773] = spike773;        spike_register[774] = spike774;        spike_register[775] = spike775;        spike_register[776] = spike776;        spike_register[777] = spike777;        spike_register[778] = spike778;        spike_register[779] = spike779;        spike_register[780] = spike780;        spike_register[781] = spike781;        spike_register[782] = spike782;        spike_register[783] = spike783;        spike_register[784] = spike784;        spike_register[785] = spike785;        spike_register[786] = spike786;        spike_register[787] = spike787;        spike_register[788] = spike788;        spike_register[789] = spike789;        spike_register[790] = spike790;        spike_register[791] = spike791;        spike_register[792] = spike792;        spike_register[793] = spike793;        spike_register[794] = spike794;        spike_register[795] = spike795;        spike_register[796] = spike796;        spike_register[797] = spike797;        spike_register[798] = spike798;        spike_register[799] = spike799;
        #0.5
        if(clear == 1'b0) begin
            for(i16 = 750; i16 <=799; i16= i16+1) begin
                if(spike_register[i16] == 1 && lock16 == 0) begin
                    lock16 = 1;
                    for(j16 = connection_pointer[i16]; j16 < connection_pointer[i16+1]; j16= j16+1) begin
                        packet16 = #0.1 {neuron_addresses[i16], downstream_connections[j16]};
                    end
                    spike_register[i16] = 0;
                    lock16 = 0;
                end
            end
        end

    end
    always @(clear, lock17, spike800, spike801, spike802, spike803, spike804, spike805, spike806, spike807, spike808, spike809, spike810, spike811, spike812, spike813, spike814, spike815, spike816, spike817, spike818, spike819, spike820, spike821, spike822, spike823, spike824, spike825, spike826, spike827, spike828, spike829, spike830, spike831, spike832, spike833, spike834, spike835, spike836, spike837, spike838, spike839, spike840, spike841, spike842, spike843, spike844, spike845, spike846, spike847, spike848, spike849) begin
        spike_register[800] = spike800;

        spike_register[801] = spike801;        spike_register[802] = spike802;        spike_register[803] = spike803;        spike_register[804] = spike804;        spike_register[805] = spike805;        spike_register[806] = spike806;        spike_register[807] = spike807;        spike_register[808] = spike808;        spike_register[809] = spike809;        spike_register[810] = spike810;        spike_register[811] = spike811;        spike_register[812] = spike812;        spike_register[813] = spike813;        spike_register[814] = spike814;        spike_register[815] = spike815;        spike_register[816] = spike816;        spike_register[817] = spike817;        spike_register[818] = spike818;        spike_register[819] = spike819;        spike_register[820] = spike820;        spike_register[821] = spike821;        spike_register[822] = spike822;        spike_register[823] = spike823;        spike_register[824] = spike824;        spike_register[825] = spike825;        spike_register[826] = spike826;        spike_register[827] = spike827;        spike_register[828] = spike828;        spike_register[829] = spike829;        spike_register[830] = spike830;        spike_register[831] = spike831;        spike_register[832] = spike832;        spike_register[833] = spike833;        spike_register[834] = spike834;        spike_register[835] = spike835;        spike_register[836] = spike836;        spike_register[837] = spike837;        spike_register[838] = spike838;        spike_register[839] = spike839;        spike_register[840] = spike840;        spike_register[841] = spike841;        spike_register[842] = spike842;        spike_register[843] = spike843;        spike_register[844] = spike844;        spike_register[845] = spike845;        spike_register[846] = spike846;        spike_register[847] = spike847;        spike_register[848] = spike848;        spike_register[849] = spike849;
        #0.5
        if(clear == 1'b0) begin
            for(i17 = 800; i17 <=849; i17= i17+1) begin
                if(spike_register[i17] == 1 && lock17 == 0) begin
                    lock17 = 1;
                    for(j17 = connection_pointer[i17]; j17 < connection_pointer[i17+1]; j17= j17+1) begin
                        packet17 = #0.1 {neuron_addresses[i17], downstream_connections[j17]};
                    end
                    spike_register[i17] = 0;
                    lock17 = 0;
                end
            end
        end

    end
    always @(clear, lock18, spike850, spike851, spike852, spike853, spike854, spike855, spike856, spike857, spike858, spike859, spike860, spike861, spike862, spike863, spike864, spike865, spike866, spike867, spike868, spike869, spike870, spike871, spike872, spike873, spike874, spike875, spike876, spike877, spike878, spike879, spike880, spike881, spike882, spike883, spike884, spike885, spike886, spike887, spike888, spike889, spike890, spike891, spike892, spike893, spike894, spike895, spike896, spike897, spike898, spike899) begin
        spike_register[850] = spike850;        spike_register[851] = spike851;        spike_register[852] = spike852;        spike_register[853] = spike853;        spike_register[854] = spike854;        spike_register[855] = spike855;        spike_register[856] = spike856;        spike_register[857] = spike857;        spike_register[858] = spike858;        spike_register[859] = spike859;        spike_register[860] = spike860;        spike_register[861] = spike861;        spike_register[862] = spike862;        spike_register[863] = spike863;        spike_register[864] = spike864;        spike_register[865] = spike865;        spike_register[866] = spike866;        spike_register[867] = spike867;        spike_register[868] = spike868;        spike_register[869] = spike869;        spike_register[870] = spike870;        spike_register[871] = spike871;        spike_register[872] = spike872;        spike_register[873] = spike873;        spike_register[874] = spike874;        spike_register[875] = spike875;        spike_register[876] = spike876;        spike_register[877] = spike877;        spike_register[878] = spike878;        spike_register[879] = spike879;        spike_register[880] = spike880;        spike_register[881] = spike881;        spike_register[882] = spike882;        spike_register[883] = spike883;        spike_register[884] = spike884;        spike_register[885] = spike885;        spike_register[886] = spike886;        spike_register[887] = spike887;        spike_register[888] = spike888;        spike_register[889] = spike889;        spike_register[890] = spike890;        spike_register[891] = spike891;        spike_register[892] = spike892;        spike_register[893] = spike893;        spike_register[894] = spike894;        spike_register[895] = spike895;        spike_register[896] = spike896;        spike_register[897] = spike897;        spike_register[898] = spike898;        spike_register[899] = spike899;
        #0.5
        if(clear == 1'b0) begin
            for(i18 = 850; i18 <=899; i18= i18+1) begin
                if(spike_register[i18] == 1 && lock18 == 0) begin
                    lock18 = 1;
                    for(j18 = connection_pointer[i18]; j18 < connection_pointer[i18+1]; j18= j18+1) begin
                        packet18 = #0.1 {neuron_addresses[i18], downstream_connections[j18]};
                    end
                    spike_register[i18] = 0;
                    lock18 = 0;
                end
            end
        end

    end
    always @(clear, lock19, spike900, spike901, spike902, spike903, spike904, spike905, spike906, spike907, spike908, spike909, spike910, spike911, spike912, spike913, spike914, spike915, spike916, spike917, spike918, spike919, spike920, spike921, spike922, spike923, spike924, spike925, spike926, spike927, spike928, spike929, spike930, spike931, spike932, spike933, spike934, spike935, spike936, spike937, spike938, spike939, spike940, spike941, spike942, spike943, spike944, spike945, spike946, spike947, spike948, spike949) begin
        spike_register[900] = spike900;

        spike_register[901] = spike901;        spike_register[902] = spike902;        spike_register[903] = spike903;        spike_register[904] = spike904;        spike_register[905] = spike905;        spike_register[906] = spike906;        spike_register[907] = spike907;        spike_register[908] = spike908;        spike_register[909] = spike909;        spike_register[910] = spike910;        spike_register[911] = spike911;        spike_register[912] = spike912;        spike_register[913] = spike913;        spike_register[914] = spike914;        spike_register[915] = spike915;        spike_register[916] = spike916;        spike_register[917] = spike917;        spike_register[918] = spike918;        spike_register[919] = spike919;        spike_register[920] = spike920;        spike_register[921] = spike921;        spike_register[922] = spike922;        spike_register[923] = spike923;        spike_register[924] = spike924;        spike_register[925] = spike925;        spike_register[926] = spike926;        spike_register[927] = spike927;        spike_register[928] = spike928;        spike_register[929] = spike929;        spike_register[930] = spike930;        spike_register[931] = spike931;        spike_register[932] = spike932;        spike_register[933] = spike933;        spike_register[934] = spike934;        spike_register[935] = spike935;        spike_register[936] = spike936;        spike_register[937] = spike937;        spike_register[938] = spike938;        spike_register[939] = spike939;        spike_register[940] = spike940;        spike_register[941] = spike941;        spike_register[942] = spike942;        spike_register[943] = spike943;        spike_register[944] = spike944;        spike_register[945] = spike945;        spike_register[946] = spike946;        spike_register[947] = spike947;        spike_register[948] = spike948;        spike_register[949] = spike949;
        #0.5
        if(clear == 1'b0) begin
            for(i19 = 900; i19 <=949; i19= i19+1) begin
                if(spike_register[i19] == 1 && lock19 == 0) begin
                    lock19 = 1;
                    for(j19 = connection_pointer[i19]; j19 < connection_pointer[i19+1]; j19= j19+1) begin
                        packet19 = #0.1 {neuron_addresses[i19], downstream_connections[j19]};
                    end
                    spike_register[i19] = 0;
                    lock19 = 0;
                end
            end
        end

    end
    always @(clear, lock20, spike950, spike951, spike952, spike953, spike954, spike955, spike956, spike957, spike958, spike959, spike960, spike961, spike962, spike963, spike964, spike965, spike966, spike967, spike968, spike969, spike970, spike971, spike972, spike973, spike974, spike975, spike976, spike977, spike978, spike979, spike980, spike981, spike982, spike983, spike984, spike985, spike986, spike987, spike988, spike989, spike990, spike991, spike992, spike993, spike994, spike995, spike996, spike997, spike998, spike999) begin
        spike_register[950] = spike950;        spike_register[951] = spike951;        spike_register[952] = spike952;        spike_register[953] = spike953;        spike_register[954] = spike954;        spike_register[955] = spike955;        spike_register[956] = spike956;        spike_register[957] = spike957;        spike_register[958] = spike958;        spike_register[959] = spike959;        spike_register[960] = spike960;        spike_register[961] = spike961;        spike_register[962] = spike962;        spike_register[963] = spike963;        spike_register[964] = spike964;        spike_register[965] = spike965;        spike_register[966] = spike966;        spike_register[967] = spike967;        spike_register[968] = spike968;        spike_register[969] = spike969;        spike_register[970] = spike970;        spike_register[971] = spike971;        spike_register[972] = spike972;        spike_register[973] = spike973;        spike_register[974] = spike974;        spike_register[975] = spike975;        spike_register[976] = spike976;        spike_register[977] = spike977;        spike_register[978] = spike978;        spike_register[979] = spike979;        spike_register[980] = spike980;        spike_register[981] = spike981;        spike_register[982] = spike982;        spike_register[983] = spike983;        spike_register[984] = spike984;        spike_register[985] = spike985;        spike_register[986] = spike986;        spike_register[987] = spike987;        spike_register[988] = spike988;        spike_register[989] = spike989;        spike_register[990] = spike990;        spike_register[991] = spike991;        spike_register[992] = spike992;        spike_register[993] = spike993;        spike_register[994] = spike994;        spike_register[995] = spike995;        spike_register[996] = spike996;        spike_register[997] = spike997;        spike_register[998] = spike998;        spike_register[999] = spike999;
        #0.5
        if(clear == 1'b0) begin
            for(i20 = 950; i20 <=999; i20= i20+1) begin
                if(spike_register[i20] == 1 && lock20 == 0) begin
                    lock20 = 1;
                    for(j20 = connection_pointer[i20]; j20 < connection_pointer[i20+1]; j20= j20+1) begin
                        packet20 = #0.1 {neuron_addresses[i20], downstream_connections[j20]};
                    end
                    spike_register[i20] = 0;
                    lock20 = 0;
                end
            end
        end

    end
    always @(clear, lock21, spike1000, spike1001, spike1002, spike1003, spike1004, spike1005, spike1006, spike1007, spike1008, spike1009, spike1010, spike1011, spike1012, spike1013, spike1014, spike1015, spike1016, spike1017, spike1018, spike1019, spike1020, spike1021, spike1022, spike1023) begin
        spike_register[1000] = spike1000;

        spike_register[1001] = spike1001;        spike_register[1002] = spike1002;        spike_register[1003] = spike1003;        spike_register[1004] = spike1004;        spike_register[1005] = spike1005;        spike_register[1006] = spike1006;        spike_register[1007] = spike1007;        spike_register[1008] = spike1008;        spike_register[1009] = spike1009;        spike_register[1010] = spike1010;        spike_register[1011] = spike1011;        spike_register[1012] = spike1012;        spike_register[1013] = spike1013;        spike_register[1014] = spike1014;        spike_register[1015] = spike1015;        spike_register[1016] = spike1016;        spike_register[1017] = spike1017;        spike_register[1018] = spike1018;        spike_register[1019] = spike1019;        spike_register[1020] = spike1020;        spike_register[1021] = spike1021;        spike_register[1022] = spike1022;        spike_register[1023] = spike1023;
        #0.5
        if(clear == 1'b0) begin
            for(i21 = 1000; i21 <=1049; i21= i21+1) begin
                if(spike_register[i21] == 1 && lock21 == 0) begin
                    lock21 = 1;
                    for(j21 = connection_pointer[i21]; j21 < connection_pointer[i21+1]; j21= j21+1) begin
                        packet21 = #0.1 {neuron_addresses[i21], downstream_connections[j21]};
                    end
                    spike_register[i21] = 0;
                    lock21 = 0;
                end
            end
        end

    end
    always @(packet1) begin 
        spike_origin = packet1[23:12];
        spike_destination = packet1[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet2) begin 
        spike_origin = packet2[23:12];
        spike_destination = packet2[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet3) begin 
        spike_origin = packet3[23:12];
        spike_destination = packet3[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet4) begin 
        spike_origin = packet4[23:12];
        spike_destination = packet4[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet5) begin 
        spike_origin = packet5[23:12];
        spike_destination = packet5[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet6) begin 
        spike_origin = packet6[23:12];
        spike_destination = packet6[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet7) begin 
        spike_origin = packet7[23:12];
        spike_destination = packet7[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet8) begin 
        spike_origin = packet8[23:12];
        spike_destination = packet8[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet9) begin 
        spike_origin = packet9[23:12];
        spike_destination = packet9[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet10) begin 
        spike_origin = packet10[23:12];
        spike_destination = packet10[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet11) begin 
        spike_origin = packet11[23:12];
        spike_destination = packet11[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet12) begin 
        spike_origin = packet12[23:12];
        spike_destination = packet12[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet13) begin 
        spike_origin = packet13[23:12];
        spike_destination = packet13[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet14) begin 
        spike_origin = packet14[23:12];
        spike_destination = packet14[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet15) begin 
        spike_origin = packet15[23:12];
        spike_destination = packet15[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet16) begin 
        spike_origin = packet16[23:12];
        spike_destination = packet16[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet17) begin 
        spike_origin = packet17[23:12];
        spike_destination = packet17[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet18) begin 
        spike_origin = packet18[23:12];
        spike_destination = packet18[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet19) begin 
        spike_origin = packet19[23:12];
        spike_destination = packet19[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet20) begin 
        spike_origin = packet20[23:12];
        spike_destination = packet20[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(packet21) begin 
        spike_origin = packet21[23:12];
        spike_destination = packet21[11:0];
        source_addresses[spike_destination] = spike_origin;
    end
    always @(spike_out_source_array[0]) begin 
        spike_out_source0 = spike_out_source_array[0];
    end
    always @(spike_out_source_array[1]) begin 
        spike_out_source1 = spike_out_source_array[1];
    end
    always @(spike_out_source_array[2]) begin 
        spike_out_source2 = spike_out_source_array[2];
    end
    always @(spike_out_source_array[3]) begin 
        spike_out_source3 = spike_out_source_array[3];
    end
    always @(spike_out_source_array[4]) begin 
        spike_out_source4 = spike_out_source_array[4];
    end
    always @(spike_out_source_array[5]) begin 
        spike_out_source5 = spike_out_source_array[5];
    end
    always @(spike_out_source_array[6]) begin 
        spike_out_source6 = spike_out_source_array[6];
    end
    always @(spike_out_source_array[7]) begin 
        spike_out_source7 = spike_out_source_array[7];
    end
    always @(spike_out_source_array[8]) begin 
        spike_out_source8 = spike_out_source_array[8];
    end
    always @(spike_out_source_array[9]) begin 
        spike_out_source9 = spike_out_source_array[9];
    end
    always @(spike_out_source_array[10]) begin 
        spike_out_source10 = spike_out_source_array[10];
    end
    always @(spike_out_source_array[11]) begin 
        spike_out_source11 = spike_out_source_array[11];
    end
    always @(spike_out_source_array[12]) begin 
        spike_out_source12 = spike_out_source_array[12];
    end
    always @(spike_out_source_array[13]) begin 
        spike_out_source13 = spike_out_source_array[13];
    end
    always @(spike_out_source_array[14]) begin 
        spike_out_source14 = spike_out_source_array[14];
    end
    always @(spike_out_source_array[15]) begin 
        spike_out_source15 = spike_out_source_array[15];
    end
    always @(spike_out_source_array[16]) begin 
        spike_out_source16 = spike_out_source_array[16];
    end
    always @(spike_out_source_array[17]) begin 
        spike_out_source17 = spike_out_source_array[17];
    end
    always @(spike_out_source_array[18]) begin 
        spike_out_source18 = spike_out_source_array[18];
    end
    always @(spike_out_source_array[19]) begin 
        spike_out_source19 = spike_out_source_array[19];
    end
    always @(spike_out_source_array[20]) begin 
        spike_out_source20 = spike_out_source_array[20];
    end
    always @(spike_out_source_array[21]) begin 
        spike_out_source21 = spike_out_source_array[21];
    end
    always @(spike_out_source_array[22]) begin 
        spike_out_source22 = spike_out_source_array[22];
    end
    always @(spike_out_source_array[23]) begin 
        spike_out_source23 = spike_out_source_array[23];
    end
    always @(spike_out_source_array[24]) begin 
        spike_out_source24 = spike_out_source_array[24];
    end
    always @(spike_out_source_array[25]) begin 
        spike_out_source25 = spike_out_source_array[25];
    end
    always @(spike_out_source_array[26]) begin 
        spike_out_source26 = spike_out_source_array[26];
    end
    always @(spike_out_source_array[27]) begin 
        spike_out_source27 = spike_out_source_array[27];
    end
    always @(spike_out_source_array[28]) begin 
        spike_out_source28 = spike_out_source_array[28];
    end
    always @(spike_out_source_array[29]) begin 
        spike_out_source29 = spike_out_source_array[29];
    end
    always @(spike_out_source_array[30]) begin 
        spike_out_source30 = spike_out_source_array[30];
    end
    always @(spike_out_source_array[31]) begin 
        spike_out_source31 = spike_out_source_array[31];
    end
    always @(spike_out_source_array[32]) begin 
        spike_out_source32 = spike_out_source_array[32];
    end
    always @(spike_out_source_array[33]) begin 
        spike_out_source33 = spike_out_source_array[33];
    end
    always @(spike_out_source_array[34]) begin 
        spike_out_source34 = spike_out_source_array[34];
    end
    always @(spike_out_source_array[35]) begin 
        spike_out_source35 = spike_out_source_array[35];
    end
    always @(spike_out_source_array[36]) begin 
        spike_out_source36 = spike_out_source_array[36];
    end
    always @(spike_out_source_array[37]) begin 
        spike_out_source37 = spike_out_source_array[37];
    end
    always @(spike_out_source_array[38]) begin 
        spike_out_source38 = spike_out_source_array[38];
    end
    always @(spike_out_source_array[39]) begin 
        spike_out_source39 = spike_out_source_array[39];
    end
    always @(spike_out_source_array[40]) begin 
        spike_out_source40 = spike_out_source_array[40];
    end
    always @(spike_out_source_array[41]) begin 
        spike_out_source41 = spike_out_source_array[41];
    end
    always @(spike_out_source_array[42]) begin 
        spike_out_source42 = spike_out_source_array[42];
    end
    always @(spike_out_source_array[43]) begin 
        spike_out_source43 = spike_out_source_array[43];
    end
    always @(spike_out_source_array[44]) begin 
        spike_out_source44 = spike_out_source_array[44];
    end
    always @(spike_out_source_array[45]) begin 
        spike_out_source45 = spike_out_source_array[45];
    end
    always @(spike_out_source_array[46]) begin 
        spike_out_source46 = spike_out_source_array[46];
    end
    always @(spike_out_source_array[47]) begin 
        spike_out_source47 = spike_out_source_array[47];
    end
    always @(spike_out_source_array[48]) begin 
        spike_out_source48 = spike_out_source_array[48];
    end
    always @(spike_out_source_array[49]) begin 
        spike_out_source49 = spike_out_source_array[49];
    end
    always @(spike_out_source_array[50]) begin 
        spike_out_source50 = spike_out_source_array[50];
    end
    always @(spike_out_source_array[51]) begin 
        spike_out_source51 = spike_out_source_array[51];
    end
    always @(spike_out_source_array[52]) begin 
        spike_out_source52 = spike_out_source_array[52];
    end
    always @(spike_out_source_array[53]) begin 
        spike_out_source53 = spike_out_source_array[53];
    end
    always @(spike_out_source_array[54]) begin 
        spike_out_source54 = spike_out_source_array[54];
    end
    always @(spike_out_source_array[55]) begin 
        spike_out_source55 = spike_out_source_array[55];
    end
    always @(spike_out_source_array[56]) begin 
        spike_out_source56 = spike_out_source_array[56];
    end
    always @(spike_out_source_array[57]) begin 
        spike_out_source57 = spike_out_source_array[57];
    end
    always @(spike_out_source_array[58]) begin 
        spike_out_source58 = spike_out_source_array[58];
    end
    always @(spike_out_source_array[59]) begin 
        spike_out_source59 = spike_out_source_array[59];
    end
    always @(spike_out_source_array[60]) begin 
        spike_out_source60 = spike_out_source_array[60];
    end
    always @(spike_out_source_array[61]) begin 
        spike_out_source61 = spike_out_source_array[61];
    end
    always @(spike_out_source_array[62]) begin 
        spike_out_source62 = spike_out_source_array[62];
    end
    always @(spike_out_source_array[63]) begin 
        spike_out_source63 = spike_out_source_array[63];
    end
    always @(spike_out_source_array[64]) begin 
        spike_out_source64 = spike_out_source_array[64];
    end
    always @(spike_out_source_array[65]) begin 
        spike_out_source65 = spike_out_source_array[65];
    end
    always @(spike_out_source_array[66]) begin 
        spike_out_source66 = spike_out_source_array[66];
    end
    always @(spike_out_source_array[67]) begin 
        spike_out_source67 = spike_out_source_array[67];
    end
    always @(spike_out_source_array[68]) begin 
        spike_out_source68 = spike_out_source_array[68];
    end
    always @(spike_out_source_array[69]) begin 
        spike_out_source69 = spike_out_source_array[69];
    end
    always @(spike_out_source_array[70]) begin 
        spike_out_source70 = spike_out_source_array[70];
    end
    always @(spike_out_source_array[71]) begin 
        spike_out_source71 = spike_out_source_array[71];
    end
    always @(spike_out_source_array[72]) begin 
        spike_out_source72 = spike_out_source_array[72];
    end
    always @(spike_out_source_array[73]) begin 
        spike_out_source73 = spike_out_source_array[73];
    end
    always @(spike_out_source_array[74]) begin 
        spike_out_source74 = spike_out_source_array[74];
    end
    always @(spike_out_source_array[75]) begin 
        spike_out_source75 = spike_out_source_array[75];
    end
    always @(spike_out_source_array[76]) begin 
        spike_out_source76 = spike_out_source_array[76];
    end
    always @(spike_out_source_array[77]) begin 
        spike_out_source77 = spike_out_source_array[77];
    end
    always @(spike_out_source_array[78]) begin 
        spike_out_source78 = spike_out_source_array[78];
    end
    always @(spike_out_source_array[79]) begin 
        spike_out_source79 = spike_out_source_array[79];
    end
    always @(spike_out_source_array[80]) begin 
        spike_out_source80 = spike_out_source_array[80];
    end
    always @(spike_out_source_array[81]) begin 
        spike_out_source81 = spike_out_source_array[81];
    end
    always @(spike_out_source_array[82]) begin 
        spike_out_source82 = spike_out_source_array[82];
    end
    always @(spike_out_source_array[83]) begin 
        spike_out_source83 = spike_out_source_array[83];
    end
    always @(spike_out_source_array[84]) begin 
        spike_out_source84 = spike_out_source_array[84];
    end
    always @(spike_out_source_array[85]) begin 
        spike_out_source85 = spike_out_source_array[85];
    end
    always @(spike_out_source_array[86]) begin 
        spike_out_source86 = spike_out_source_array[86];
    end
    always @(spike_out_source_array[87]) begin 
        spike_out_source87 = spike_out_source_array[87];
    end
    always @(spike_out_source_array[88]) begin 
        spike_out_source88 = spike_out_source_array[88];
    end
    always @(spike_out_source_array[89]) begin 
        spike_out_source89 = spike_out_source_array[89];
    end
    always @(spike_out_source_array[90]) begin 
        spike_out_source90 = spike_out_source_array[90];
    end
    always @(spike_out_source_array[91]) begin 
        spike_out_source91 = spike_out_source_array[91];
    end
    always @(spike_out_source_array[92]) begin 
        spike_out_source92 = spike_out_source_array[92];
    end
    always @(spike_out_source_array[93]) begin 
        spike_out_source93 = spike_out_source_array[93];
    end
    always @(spike_out_source_array[94]) begin 
        spike_out_source94 = spike_out_source_array[94];
    end
    always @(spike_out_source_array[95]) begin 
        spike_out_source95 = spike_out_source_array[95];
    end
    always @(spike_out_source_array[96]) begin 
        spike_out_source96 = spike_out_source_array[96];
    end
    always @(spike_out_source_array[97]) begin 
        spike_out_source97 = spike_out_source_array[97];
    end
    always @(spike_out_source_array[98]) begin 
        spike_out_source98 = spike_out_source_array[98];
    end
    always @(spike_out_source_array[99]) begin 
        spike_out_source99 = spike_out_source_array[99];
    end
    always @(spike_out_source_array[100]) begin 
        spike_out_source100 = spike_out_source_array[100];
    end
    always @(spike_out_source_array[101]) begin 
        spike_out_source101 = spike_out_source_array[101];
    end
    always @(spike_out_source_array[102]) begin 
        spike_out_source102 = spike_out_source_array[102];
    end
    always @(spike_out_source_array[103]) begin 
        spike_out_source103 = spike_out_source_array[103];
    end
    always @(spike_out_source_array[104]) begin 
        spike_out_source104 = spike_out_source_array[104];
    end
    always @(spike_out_source_array[105]) begin 
        spike_out_source105 = spike_out_source_array[105];
    end
    always @(spike_out_source_array[106]) begin 
        spike_out_source106 = spike_out_source_array[106];
    end
    always @(spike_out_source_array[107]) begin 
        spike_out_source107 = spike_out_source_array[107];
    end
    always @(spike_out_source_array[108]) begin 
        spike_out_source108 = spike_out_source_array[108];
    end
    always @(spike_out_source_array[109]) begin 
        spike_out_source109 = spike_out_source_array[109];
    end
    always @(spike_out_source_array[110]) begin 
        spike_out_source110 = spike_out_source_array[110];
    end
    always @(spike_out_source_array[111]) begin 
        spike_out_source111 = spike_out_source_array[111];
    end
    always @(spike_out_source_array[112]) begin 
        spike_out_source112 = spike_out_source_array[112];
    end
    always @(spike_out_source_array[113]) begin 
        spike_out_source113 = spike_out_source_array[113];
    end
    always @(spike_out_source_array[114]) begin 
        spike_out_source114 = spike_out_source_array[114];
    end
    always @(spike_out_source_array[115]) begin 
        spike_out_source115 = spike_out_source_array[115];
    end
    always @(spike_out_source_array[116]) begin 
        spike_out_source116 = spike_out_source_array[116];
    end
    always @(spike_out_source_array[117]) begin 
        spike_out_source117 = spike_out_source_array[117];
    end
    always @(spike_out_source_array[118]) begin 
        spike_out_source118 = spike_out_source_array[118];
    end
    always @(spike_out_source_array[119]) begin 
        spike_out_source119 = spike_out_source_array[119];
    end
    always @(spike_out_source_array[120]) begin 
        spike_out_source120 = spike_out_source_array[120];
    end
    always @(spike_out_source_array[121]) begin 
        spike_out_source121 = spike_out_source_array[121];
    end
    always @(spike_out_source_array[122]) begin 
        spike_out_source122 = spike_out_source_array[122];
    end
    always @(spike_out_source_array[123]) begin 
        spike_out_source123 = spike_out_source_array[123];
    end
    always @(spike_out_source_array[124]) begin 
        spike_out_source124 = spike_out_source_array[124];
    end
    always @(spike_out_source_array[125]) begin 
        spike_out_source125 = spike_out_source_array[125];
    end
    always @(spike_out_source_array[126]) begin 
        spike_out_source126 = spike_out_source_array[126];
    end
    always @(spike_out_source_array[127]) begin 
        spike_out_source127 = spike_out_source_array[127];
    end
    always @(spike_out_source_array[128]) begin 
        spike_out_source128 = spike_out_source_array[128];
    end
    always @(spike_out_source_array[129]) begin 
        spike_out_source129 = spike_out_source_array[129];
    end
    always @(spike_out_source_array[130]) begin 
        spike_out_source130 = spike_out_source_array[130];
    end
    always @(spike_out_source_array[131]) begin 
        spike_out_source131 = spike_out_source_array[131];
    end
    always @(spike_out_source_array[132]) begin 
        spike_out_source132 = spike_out_source_array[132];
    end
    always @(spike_out_source_array[133]) begin 
        spike_out_source133 = spike_out_source_array[133];
    end
    always @(spike_out_source_array[134]) begin 
        spike_out_source134 = spike_out_source_array[134];
    end
    always @(spike_out_source_array[135]) begin 
        spike_out_source135 = spike_out_source_array[135];
    end
    always @(spike_out_source_array[136]) begin 
        spike_out_source136 = spike_out_source_array[136];
    end
    always @(spike_out_source_array[137]) begin 
        spike_out_source137 = spike_out_source_array[137];
    end
    always @(spike_out_source_array[138]) begin 
        spike_out_source138 = spike_out_source_array[138];
    end
    always @(spike_out_source_array[139]) begin 
        spike_out_source139 = spike_out_source_array[139];
    end
    always @(spike_out_source_array[140]) begin 
        spike_out_source140 = spike_out_source_array[140];
    end
    always @(spike_out_source_array[141]) begin 
        spike_out_source141 = spike_out_source_array[141];
    end
    always @(spike_out_source_array[142]) begin 
        spike_out_source142 = spike_out_source_array[142];
    end
    always @(spike_out_source_array[143]) begin 
        spike_out_source143 = spike_out_source_array[143];
    end
    always @(spike_out_source_array[144]) begin 
        spike_out_source144 = spike_out_source_array[144];
    end
    always @(spike_out_source_array[145]) begin 
        spike_out_source145 = spike_out_source_array[145];
    end
    always @(spike_out_source_array[146]) begin 
        spike_out_source146 = spike_out_source_array[146];
    end
    always @(spike_out_source_array[147]) begin 
        spike_out_source147 = spike_out_source_array[147];
    end
    always @(spike_out_source_array[148]) begin 
        spike_out_source148 = spike_out_source_array[148];
    end
    always @(spike_out_source_array[149]) begin 
        spike_out_source149 = spike_out_source_array[149];
    end
    always @(spike_out_source_array[150]) begin 
        spike_out_source150 = spike_out_source_array[150];
    end
    always @(spike_out_source_array[151]) begin 
        spike_out_source151 = spike_out_source_array[151];
    end
    always @(spike_out_source_array[152]) begin 
        spike_out_source152 = spike_out_source_array[152];
    end
    always @(spike_out_source_array[153]) begin 
        spike_out_source153 = spike_out_source_array[153];
    end
    always @(spike_out_source_array[154]) begin 
        spike_out_source154 = spike_out_source_array[154];
    end
    always @(spike_out_source_array[155]) begin 
        spike_out_source155 = spike_out_source_array[155];
    end
    always @(spike_out_source_array[156]) begin 
        spike_out_source156 = spike_out_source_array[156];
    end
    always @(spike_out_source_array[157]) begin 
        spike_out_source157 = spike_out_source_array[157];
    end
    always @(spike_out_source_array[158]) begin 
        spike_out_source158 = spike_out_source_array[158];
    end
    always @(spike_out_source_array[159]) begin 
        spike_out_source159 = spike_out_source_array[159];
    end
    always @(spike_out_source_array[160]) begin 
        spike_out_source160 = spike_out_source_array[160];
    end
    always @(spike_out_source_array[161]) begin 
        spike_out_source161 = spike_out_source_array[161];
    end
    always @(spike_out_source_array[162]) begin 
        spike_out_source162 = spike_out_source_array[162];
    end
    always @(spike_out_source_array[163]) begin 
        spike_out_source163 = spike_out_source_array[163];
    end
    always @(spike_out_source_array[164]) begin 
        spike_out_source164 = spike_out_source_array[164];
    end
    always @(spike_out_source_array[165]) begin 
        spike_out_source165 = spike_out_source_array[165];
    end
    always @(spike_out_source_array[166]) begin 
        spike_out_source166 = spike_out_source_array[166];
    end
    always @(spike_out_source_array[167]) begin 
        spike_out_source167 = spike_out_source_array[167];
    end
    always @(spike_out_source_array[168]) begin 
        spike_out_source168 = spike_out_source_array[168];
    end
    always @(spike_out_source_array[169]) begin 
        spike_out_source169 = spike_out_source_array[169];
    end
    always @(spike_out_source_array[170]) begin 
        spike_out_source170 = spike_out_source_array[170];
    end
    always @(spike_out_source_array[171]) begin 
        spike_out_source171 = spike_out_source_array[171];
    end
    always @(spike_out_source_array[172]) begin 
        spike_out_source172 = spike_out_source_array[172];
    end
    always @(spike_out_source_array[173]) begin 
        spike_out_source173 = spike_out_source_array[173];
    end
    always @(spike_out_source_array[174]) begin 
        spike_out_source174 = spike_out_source_array[174];
    end
    always @(spike_out_source_array[175]) begin 
        spike_out_source175 = spike_out_source_array[175];
    end
    always @(spike_out_source_array[176]) begin 
        spike_out_source176 = spike_out_source_array[176];
    end
    always @(spike_out_source_array[177]) begin 
        spike_out_source177 = spike_out_source_array[177];
    end
    always @(spike_out_source_array[178]) begin 
        spike_out_source178 = spike_out_source_array[178];
    end
    always @(spike_out_source_array[179]) begin 
        spike_out_source179 = spike_out_source_array[179];
    end
    always @(spike_out_source_array[180]) begin 
        spike_out_source180 = spike_out_source_array[180];
    end
    always @(spike_out_source_array[181]) begin 
        spike_out_source181 = spike_out_source_array[181];
    end
    always @(spike_out_source_array[182]) begin 
        spike_out_source182 = spike_out_source_array[182];
    end
    always @(spike_out_source_array[183]) begin 
        spike_out_source183 = spike_out_source_array[183];
    end
    always @(spike_out_source_array[184]) begin 
        spike_out_source184 = spike_out_source_array[184];
    end
    always @(spike_out_source_array[185]) begin 
        spike_out_source185 = spike_out_source_array[185];
    end
    always @(spike_out_source_array[186]) begin 
        spike_out_source186 = spike_out_source_array[186];
    end
    always @(spike_out_source_array[187]) begin 
        spike_out_source187 = spike_out_source_array[187];
    end
    always @(spike_out_source_array[188]) begin 
        spike_out_source188 = spike_out_source_array[188];
    end
    always @(spike_out_source_array[189]) begin 
        spike_out_source189 = spike_out_source_array[189];
    end
    always @(spike_out_source_array[190]) begin 
        spike_out_source190 = spike_out_source_array[190];
    end
    always @(spike_out_source_array[191]) begin 
        spike_out_source191 = spike_out_source_array[191];
    end
    always @(spike_out_source_array[192]) begin 
        spike_out_source192 = spike_out_source_array[192];
    end
    always @(spike_out_source_array[193]) begin 
        spike_out_source193 = spike_out_source_array[193];
    end
    always @(spike_out_source_array[194]) begin 
        spike_out_source194 = spike_out_source_array[194];
    end
    always @(spike_out_source_array[195]) begin 
        spike_out_source195 = spike_out_source_array[195];
    end
    always @(spike_out_source_array[196]) begin 
        spike_out_source196 = spike_out_source_array[196];
    end
    always @(spike_out_source_array[197]) begin 
        spike_out_source197 = spike_out_source_array[197];
    end
    always @(spike_out_source_array[198]) begin 
        spike_out_source198 = spike_out_source_array[198];
    end
    always @(spike_out_source_array[199]) begin 
        spike_out_source199 = spike_out_source_array[199];
    end
    always @(spike_out_source_array[200]) begin 
        spike_out_source200 = spike_out_source_array[200];
    end
    always @(spike_out_source_array[201]) begin 
        spike_out_source201 = spike_out_source_array[201];
    end
    always @(spike_out_source_array[202]) begin 
        spike_out_source202 = spike_out_source_array[202];
    end
    always @(spike_out_source_array[203]) begin 
        spike_out_source203 = spike_out_source_array[203];
    end
    always @(spike_out_source_array[204]) begin 
        spike_out_source204 = spike_out_source_array[204];
    end
    always @(spike_out_source_array[205]) begin 
        spike_out_source205 = spike_out_source_array[205];
    end
    always @(spike_out_source_array[206]) begin 
        spike_out_source206 = spike_out_source_array[206];
    end
    always @(spike_out_source_array[207]) begin 
        spike_out_source207 = spike_out_source_array[207];
    end
    always @(spike_out_source_array[208]) begin 
        spike_out_source208 = spike_out_source_array[208];
    end
    always @(spike_out_source_array[209]) begin 
        spike_out_source209 = spike_out_source_array[209];
    end
    always @(spike_out_source_array[210]) begin 
        spike_out_source210 = spike_out_source_array[210];
    end
    always @(spike_out_source_array[211]) begin 
        spike_out_source211 = spike_out_source_array[211];
    end
    always @(spike_out_source_array[212]) begin 
        spike_out_source212 = spike_out_source_array[212];
    end
    always @(spike_out_source_array[213]) begin 
        spike_out_source213 = spike_out_source_array[213];
    end
    always @(spike_out_source_array[214]) begin 
        spike_out_source214 = spike_out_source_array[214];
    end
    always @(spike_out_source_array[215]) begin 
        spike_out_source215 = spike_out_source_array[215];
    end
    always @(spike_out_source_array[216]) begin 
        spike_out_source216 = spike_out_source_array[216];
    end
    always @(spike_out_source_array[217]) begin 
        spike_out_source217 = spike_out_source_array[217];
    end
    always @(spike_out_source_array[218]) begin 
        spike_out_source218 = spike_out_source_array[218];
    end
    always @(spike_out_source_array[219]) begin 
        spike_out_source219 = spike_out_source_array[219];
    end
    always @(spike_out_source_array[220]) begin 
        spike_out_source220 = spike_out_source_array[220];
    end
    always @(spike_out_source_array[221]) begin 
        spike_out_source221 = spike_out_source_array[221];
    end
    always @(spike_out_source_array[222]) begin 
        spike_out_source222 = spike_out_source_array[222];
    end
    always @(spike_out_source_array[223]) begin 
        spike_out_source223 = spike_out_source_array[223];
    end
    always @(spike_out_source_array[224]) begin 
        spike_out_source224 = spike_out_source_array[224];
    end
    always @(spike_out_source_array[225]) begin 
        spike_out_source225 = spike_out_source_array[225];
    end
    always @(spike_out_source_array[226]) begin 
        spike_out_source226 = spike_out_source_array[226];
    end
    always @(spike_out_source_array[227]) begin 
        spike_out_source227 = spike_out_source_array[227];
    end
    always @(spike_out_source_array[228]) begin 
        spike_out_source228 = spike_out_source_array[228];
    end
    always @(spike_out_source_array[229]) begin 
        spike_out_source229 = spike_out_source_array[229];
    end
    always @(spike_out_source_array[230]) begin 
        spike_out_source230 = spike_out_source_array[230];
    end
    always @(spike_out_source_array[231]) begin 
        spike_out_source231 = spike_out_source_array[231];
    end
    always @(spike_out_source_array[232]) begin 
        spike_out_source232 = spike_out_source_array[232];
    end
    always @(spike_out_source_array[233]) begin 
        spike_out_source233 = spike_out_source_array[233];
    end
    always @(spike_out_source_array[234]) begin 
        spike_out_source234 = spike_out_source_array[234];
    end
    always @(spike_out_source_array[235]) begin 
        spike_out_source235 = spike_out_source_array[235];
    end
    always @(spike_out_source_array[236]) begin 
        spike_out_source236 = spike_out_source_array[236];
    end
    always @(spike_out_source_array[237]) begin 
        spike_out_source237 = spike_out_source_array[237];
    end
    always @(spike_out_source_array[238]) begin 
        spike_out_source238 = spike_out_source_array[238];
    end
    always @(spike_out_source_array[239]) begin 
        spike_out_source239 = spike_out_source_array[239];
    end
    always @(spike_out_source_array[240]) begin 
        spike_out_source240 = spike_out_source_array[240];
    end
    always @(spike_out_source_array[241]) begin 
        spike_out_source241 = spike_out_source_array[241];
    end
    always @(spike_out_source_array[242]) begin 
        spike_out_source242 = spike_out_source_array[242];
    end
    always @(spike_out_source_array[243]) begin 
        spike_out_source243 = spike_out_source_array[243];
    end
    always @(spike_out_source_array[244]) begin 
        spike_out_source244 = spike_out_source_array[244];
    end
    always @(spike_out_source_array[245]) begin 
        spike_out_source245 = spike_out_source_array[245];
    end
    always @(spike_out_source_array[246]) begin 
        spike_out_source246 = spike_out_source_array[246];
    end
    always @(spike_out_source_array[247]) begin 
        spike_out_source247 = spike_out_source_array[247];
    end
    always @(spike_out_source_array[248]) begin 
        spike_out_source248 = spike_out_source_array[248];
    end
    always @(spike_out_source_array[249]) begin 
        spike_out_source249 = spike_out_source_array[249];
    end
    always @(spike_out_source_array[250]) begin 
        spike_out_source250 = spike_out_source_array[250];
    end
    always @(spike_out_source_array[251]) begin 
        spike_out_source251 = spike_out_source_array[251];
    end
    always @(spike_out_source_array[252]) begin 
        spike_out_source252 = spike_out_source_array[252];
    end
    always @(spike_out_source_array[253]) begin 
        spike_out_source253 = spike_out_source_array[253];
    end
    always @(spike_out_source_array[254]) begin 
        spike_out_source254 = spike_out_source_array[254];
    end
    always @(spike_out_source_array[255]) begin 
        spike_out_source255 = spike_out_source_array[255];
    end
    always @(spike_out_source_array[256]) begin 
        spike_out_source256 = spike_out_source_array[256];
    end
    always @(spike_out_source_array[257]) begin 
        spike_out_source257 = spike_out_source_array[257];
    end
    always @(spike_out_source_array[258]) begin 
        spike_out_source258 = spike_out_source_array[258];
    end
    always @(spike_out_source_array[259]) begin 
        spike_out_source259 = spike_out_source_array[259];
    end
    always @(spike_out_source_array[260]) begin 
        spike_out_source260 = spike_out_source_array[260];
    end
    always @(spike_out_source_array[261]) begin 
        spike_out_source261 = spike_out_source_array[261];
    end
    always @(spike_out_source_array[262]) begin 
        spike_out_source262 = spike_out_source_array[262];
    end
    always @(spike_out_source_array[263]) begin 
        spike_out_source263 = spike_out_source_array[263];
    end
    always @(spike_out_source_array[264]) begin 
        spike_out_source264 = spike_out_source_array[264];
    end
    always @(spike_out_source_array[265]) begin 
        spike_out_source265 = spike_out_source_array[265];
    end
    always @(spike_out_source_array[266]) begin 
        spike_out_source266 = spike_out_source_array[266];
    end
    always @(spike_out_source_array[267]) begin 
        spike_out_source267 = spike_out_source_array[267];
    end
    always @(spike_out_source_array[268]) begin 
        spike_out_source268 = spike_out_source_array[268];
    end
    always @(spike_out_source_array[269]) begin 
        spike_out_source269 = spike_out_source_array[269];
    end
    always @(spike_out_source_array[270]) begin 
        spike_out_source270 = spike_out_source_array[270];
    end
    always @(spike_out_source_array[271]) begin 
        spike_out_source271 = spike_out_source_array[271];
    end
    always @(spike_out_source_array[272]) begin 
        spike_out_source272 = spike_out_source_array[272];
    end
    always @(spike_out_source_array[273]) begin 
        spike_out_source273 = spike_out_source_array[273];
    end
    always @(spike_out_source_array[274]) begin 
        spike_out_source274 = spike_out_source_array[274];
    end
    always @(spike_out_source_array[275]) begin 
        spike_out_source275 = spike_out_source_array[275];
    end
    always @(spike_out_source_array[276]) begin 
        spike_out_source276 = spike_out_source_array[276];
    end
    always @(spike_out_source_array[277]) begin 
        spike_out_source277 = spike_out_source_array[277];
    end
    always @(spike_out_source_array[278]) begin 
        spike_out_source278 = spike_out_source_array[278];
    end
    always @(spike_out_source_array[279]) begin 
        spike_out_source279 = spike_out_source_array[279];
    end
    always @(spike_out_source_array[280]) begin 
        spike_out_source280 = spike_out_source_array[280];
    end
    always @(spike_out_source_array[281]) begin 
        spike_out_source281 = spike_out_source_array[281];
    end
    always @(spike_out_source_array[282]) begin 
        spike_out_source282 = spike_out_source_array[282];
    end
    always @(spike_out_source_array[283]) begin 
        spike_out_source283 = spike_out_source_array[283];
    end
    always @(spike_out_source_array[284]) begin 
        spike_out_source284 = spike_out_source_array[284];
    end
    always @(spike_out_source_array[285]) begin 
        spike_out_source285 = spike_out_source_array[285];
    end
    always @(spike_out_source_array[286]) begin 
        spike_out_source286 = spike_out_source_array[286];
    end
    always @(spike_out_source_array[287]) begin 
        spike_out_source287 = spike_out_source_array[287];
    end
    always @(spike_out_source_array[288]) begin 
        spike_out_source288 = spike_out_source_array[288];
    end
    always @(spike_out_source_array[289]) begin 
        spike_out_source289 = spike_out_source_array[289];
    end
    always @(spike_out_source_array[290]) begin 
        spike_out_source290 = spike_out_source_array[290];
    end
    always @(spike_out_source_array[291]) begin 
        spike_out_source291 = spike_out_source_array[291];
    end
    always @(spike_out_source_array[292]) begin 
        spike_out_source292 = spike_out_source_array[292];
    end
    always @(spike_out_source_array[293]) begin 
        spike_out_source293 = spike_out_source_array[293];
    end
    always @(spike_out_source_array[294]) begin 
        spike_out_source294 = spike_out_source_array[294];
    end
    always @(spike_out_source_array[295]) begin 
        spike_out_source295 = spike_out_source_array[295];
    end
    always @(spike_out_source_array[296]) begin 
        spike_out_source296 = spike_out_source_array[296];
    end
    always @(spike_out_source_array[297]) begin 
        spike_out_source297 = spike_out_source_array[297];
    end
    always @(spike_out_source_array[298]) begin 
        spike_out_source298 = spike_out_source_array[298];
    end
    always @(spike_out_source_array[299]) begin 
        spike_out_source299 = spike_out_source_array[299];
    end
    always @(spike_out_source_array[300]) begin 
        spike_out_source300 = spike_out_source_array[300];
    end
    always @(spike_out_source_array[301]) begin 
        spike_out_source301 = spike_out_source_array[301];
    end
    always @(spike_out_source_array[302]) begin 
        spike_out_source302 = spike_out_source_array[302];
    end
    always @(spike_out_source_array[303]) begin 
        spike_out_source303 = spike_out_source_array[303];
    end
    always @(spike_out_source_array[304]) begin 
        spike_out_source304 = spike_out_source_array[304];
    end
    always @(spike_out_source_array[305]) begin 
        spike_out_source305 = spike_out_source_array[305];
    end
    always @(spike_out_source_array[306]) begin 
        spike_out_source306 = spike_out_source_array[306];
    end
    always @(spike_out_source_array[307]) begin 
        spike_out_source307 = spike_out_source_array[307];
    end
    always @(spike_out_source_array[308]) begin 
        spike_out_source308 = spike_out_source_array[308];
    end
    always @(spike_out_source_array[309]) begin 
        spike_out_source309 = spike_out_source_array[309];
    end
    always @(spike_out_source_array[310]) begin 
        spike_out_source310 = spike_out_source_array[310];
    end
    always @(spike_out_source_array[311]) begin 
        spike_out_source311 = spike_out_source_array[311];
    end
    always @(spike_out_source_array[312]) begin 
        spike_out_source312 = spike_out_source_array[312];
    end
    always @(spike_out_source_array[313]) begin 
        spike_out_source313 = spike_out_source_array[313];
    end
    always @(spike_out_source_array[314]) begin 
        spike_out_source314 = spike_out_source_array[314];
    end
    always @(spike_out_source_array[315]) begin 
        spike_out_source315 = spike_out_source_array[315];
    end
    always @(spike_out_source_array[316]) begin 
        spike_out_source316 = spike_out_source_array[316];
    end
    always @(spike_out_source_array[317]) begin 
        spike_out_source317 = spike_out_source_array[317];
    end
    always @(spike_out_source_array[318]) begin 
        spike_out_source318 = spike_out_source_array[318];
    end
    always @(spike_out_source_array[319]) begin 
        spike_out_source319 = spike_out_source_array[319];
    end
    always @(spike_out_source_array[320]) begin 
        spike_out_source320 = spike_out_source_array[320];
    end
    always @(spike_out_source_array[321]) begin 
        spike_out_source321 = spike_out_source_array[321];
    end
    always @(spike_out_source_array[322]) begin 
        spike_out_source322 = spike_out_source_array[322];
    end
    always @(spike_out_source_array[323]) begin 
        spike_out_source323 = spike_out_source_array[323];
    end
    always @(spike_out_source_array[324]) begin 
        spike_out_source324 = spike_out_source_array[324];
    end
    always @(spike_out_source_array[325]) begin 
        spike_out_source325 = spike_out_source_array[325];
    end
    always @(spike_out_source_array[326]) begin 
        spike_out_source326 = spike_out_source_array[326];
    end
    always @(spike_out_source_array[327]) begin 
        spike_out_source327 = spike_out_source_array[327];
    end
    always @(spike_out_source_array[328]) begin 
        spike_out_source328 = spike_out_source_array[328];
    end
    always @(spike_out_source_array[329]) begin 
        spike_out_source329 = spike_out_source_array[329];
    end
    always @(spike_out_source_array[330]) begin 
        spike_out_source330 = spike_out_source_array[330];
    end
    always @(spike_out_source_array[331]) begin 
        spike_out_source331 = spike_out_source_array[331];
    end
    always @(spike_out_source_array[332]) begin 
        spike_out_source332 = spike_out_source_array[332];
    end
    always @(spike_out_source_array[333]) begin 
        spike_out_source333 = spike_out_source_array[333];
    end
    always @(spike_out_source_array[334]) begin 
        spike_out_source334 = spike_out_source_array[334];
    end
    always @(spike_out_source_array[335]) begin 
        spike_out_source335 = spike_out_source_array[335];
    end
    always @(spike_out_source_array[336]) begin 
        spike_out_source336 = spike_out_source_array[336];
    end
    always @(spike_out_source_array[337]) begin 
        spike_out_source337 = spike_out_source_array[337];
    end
    always @(spike_out_source_array[338]) begin 
        spike_out_source338 = spike_out_source_array[338];
    end
    always @(spike_out_source_array[339]) begin 
        spike_out_source339 = spike_out_source_array[339];
    end
    always @(spike_out_source_array[340]) begin 
        spike_out_source340 = spike_out_source_array[340];
    end
    always @(spike_out_source_array[341]) begin 
        spike_out_source341 = spike_out_source_array[341];
    end
    always @(spike_out_source_array[342]) begin 
        spike_out_source342 = spike_out_source_array[342];
    end
    always @(spike_out_source_array[343]) begin 
        spike_out_source343 = spike_out_source_array[343];
    end
    always @(spike_out_source_array[344]) begin 
        spike_out_source344 = spike_out_source_array[344];
    end
    always @(spike_out_source_array[345]) begin 
        spike_out_source345 = spike_out_source_array[345];
    end
    always @(spike_out_source_array[346]) begin 
        spike_out_source346 = spike_out_source_array[346];
    end
    always @(spike_out_source_array[347]) begin 
        spike_out_source347 = spike_out_source_array[347];
    end
    always @(spike_out_source_array[348]) begin 
        spike_out_source348 = spike_out_source_array[348];
    end
    always @(spike_out_source_array[349]) begin 
        spike_out_source349 = spike_out_source_array[349];
    end
    always @(spike_out_source_array[350]) begin 
        spike_out_source350 = spike_out_source_array[350];
    end
    always @(spike_out_source_array[351]) begin 
        spike_out_source351 = spike_out_source_array[351];
    end
    always @(spike_out_source_array[352]) begin 
        spike_out_source352 = spike_out_source_array[352];
    end
    always @(spike_out_source_array[353]) begin 
        spike_out_source353 = spike_out_source_array[353];
    end
    always @(spike_out_source_array[354]) begin 
        spike_out_source354 = spike_out_source_array[354];
    end
    always @(spike_out_source_array[355]) begin 
        spike_out_source355 = spike_out_source_array[355];
    end
    always @(spike_out_source_array[356]) begin 
        spike_out_source356 = spike_out_source_array[356];
    end
    always @(spike_out_source_array[357]) begin 
        spike_out_source357 = spike_out_source_array[357];
    end
    always @(spike_out_source_array[358]) begin 
        spike_out_source358 = spike_out_source_array[358];
    end
    always @(spike_out_source_array[359]) begin 
        spike_out_source359 = spike_out_source_array[359];
    end
    always @(spike_out_source_array[360]) begin 
        spike_out_source360 = spike_out_source_array[360];
    end
    always @(spike_out_source_array[361]) begin 
        spike_out_source361 = spike_out_source_array[361];
    end
    always @(spike_out_source_array[362]) begin 
        spike_out_source362 = spike_out_source_array[362];
    end
    always @(spike_out_source_array[363]) begin 
        spike_out_source363 = spike_out_source_array[363];
    end
    always @(spike_out_source_array[364]) begin 
        spike_out_source364 = spike_out_source_array[364];
    end
    always @(spike_out_source_array[365]) begin 
        spike_out_source365 = spike_out_source_array[365];
    end
    always @(spike_out_source_array[366]) begin 
        spike_out_source366 = spike_out_source_array[366];
    end
    always @(spike_out_source_array[367]) begin 
        spike_out_source367 = spike_out_source_array[367];
    end
    always @(spike_out_source_array[368]) begin 
        spike_out_source368 = spike_out_source_array[368];
    end
    always @(spike_out_source_array[369]) begin 
        spike_out_source369 = spike_out_source_array[369];
    end
    always @(spike_out_source_array[370]) begin 
        spike_out_source370 = spike_out_source_array[370];
    end
    always @(spike_out_source_array[371]) begin 
        spike_out_source371 = spike_out_source_array[371];
    end
    always @(spike_out_source_array[372]) begin 
        spike_out_source372 = spike_out_source_array[372];
    end
    always @(spike_out_source_array[373]) begin 
        spike_out_source373 = spike_out_source_array[373];
    end
    always @(spike_out_source_array[374]) begin 
        spike_out_source374 = spike_out_source_array[374];
    end
    always @(spike_out_source_array[375]) begin 
        spike_out_source375 = spike_out_source_array[375];
    end
    always @(spike_out_source_array[376]) begin 
        spike_out_source376 = spike_out_source_array[376];
    end
    always @(spike_out_source_array[377]) begin 
        spike_out_source377 = spike_out_source_array[377];
    end
    always @(spike_out_source_array[378]) begin 
        spike_out_source378 = spike_out_source_array[378];
    end
    always @(spike_out_source_array[379]) begin 
        spike_out_source379 = spike_out_source_array[379];
    end
    always @(spike_out_source_array[380]) begin 
        spike_out_source380 = spike_out_source_array[380];
    end
    always @(spike_out_source_array[381]) begin 
        spike_out_source381 = spike_out_source_array[381];
    end
    always @(spike_out_source_array[382]) begin 
        spike_out_source382 = spike_out_source_array[382];
    end
    always @(spike_out_source_array[383]) begin 
        spike_out_source383 = spike_out_source_array[383];
    end
    always @(spike_out_source_array[384]) begin 
        spike_out_source384 = spike_out_source_array[384];
    end
    always @(spike_out_source_array[385]) begin 
        spike_out_source385 = spike_out_source_array[385];
    end
    always @(spike_out_source_array[386]) begin 
        spike_out_source386 = spike_out_source_array[386];
    end
    always @(spike_out_source_array[387]) begin 
        spike_out_source387 = spike_out_source_array[387];
    end
    always @(spike_out_source_array[388]) begin 
        spike_out_source388 = spike_out_source_array[388];
    end
    always @(spike_out_source_array[389]) begin 
        spike_out_source389 = spike_out_source_array[389];
    end
    always @(spike_out_source_array[390]) begin 
        spike_out_source390 = spike_out_source_array[390];
    end
    always @(spike_out_source_array[391]) begin 
        spike_out_source391 = spike_out_source_array[391];
    end
    always @(spike_out_source_array[392]) begin 
        spike_out_source392 = spike_out_source_array[392];
    end
    always @(spike_out_source_array[393]) begin 
        spike_out_source393 = spike_out_source_array[393];
    end
    always @(spike_out_source_array[394]) begin 
        spike_out_source394 = spike_out_source_array[394];
    end
    always @(spike_out_source_array[395]) begin 
        spike_out_source395 = spike_out_source_array[395];
    end
    always @(spike_out_source_array[396]) begin 
        spike_out_source396 = spike_out_source_array[396];
    end
    always @(spike_out_source_array[397]) begin 
        spike_out_source397 = spike_out_source_array[397];
    end
    always @(spike_out_source_array[398]) begin 
        spike_out_source398 = spike_out_source_array[398];
    end
    always @(spike_out_source_array[399]) begin 
        spike_out_source399 = spike_out_source_array[399];
    end
    always @(spike_out_source_array[400]) begin 
        spike_out_source400 = spike_out_source_array[400];
    end
    always @(spike_out_source_array[401]) begin 
        spike_out_source401 = spike_out_source_array[401];
    end
    always @(spike_out_source_array[402]) begin 
        spike_out_source402 = spike_out_source_array[402];
    end
    always @(spike_out_source_array[403]) begin 
        spike_out_source403 = spike_out_source_array[403];
    end
    always @(spike_out_source_array[404]) begin 
        spike_out_source404 = spike_out_source_array[404];
    end
    always @(spike_out_source_array[405]) begin 
        spike_out_source405 = spike_out_source_array[405];
    end
    always @(spike_out_source_array[406]) begin 
        spike_out_source406 = spike_out_source_array[406];
    end
    always @(spike_out_source_array[407]) begin 
        spike_out_source407 = spike_out_source_array[407];
    end
    always @(spike_out_source_array[408]) begin 
        spike_out_source408 = spike_out_source_array[408];
    end
    always @(spike_out_source_array[409]) begin 
        spike_out_source409 = spike_out_source_array[409];
    end
    always @(spike_out_source_array[410]) begin 
        spike_out_source410 = spike_out_source_array[410];
    end
    always @(spike_out_source_array[411]) begin 
        spike_out_source411 = spike_out_source_array[411];
    end
    always @(spike_out_source_array[412]) begin 
        spike_out_source412 = spike_out_source_array[412];
    end
    always @(spike_out_source_array[413]) begin 
        spike_out_source413 = spike_out_source_array[413];
    end
    always @(spike_out_source_array[414]) begin 
        spike_out_source414 = spike_out_source_array[414];
    end
    always @(spike_out_source_array[415]) begin 
        spike_out_source415 = spike_out_source_array[415];
    end
    always @(spike_out_source_array[416]) begin 
        spike_out_source416 = spike_out_source_array[416];
    end
    always @(spike_out_source_array[417]) begin 
        spike_out_source417 = spike_out_source_array[417];
    end
    always @(spike_out_source_array[418]) begin 
        spike_out_source418 = spike_out_source_array[418];
    end
    always @(spike_out_source_array[419]) begin 
        spike_out_source419 = spike_out_source_array[419];
    end
    always @(spike_out_source_array[420]) begin 
        spike_out_source420 = spike_out_source_array[420];
    end
    always @(spike_out_source_array[421]) begin 
        spike_out_source421 = spike_out_source_array[421];
    end
    always @(spike_out_source_array[422]) begin 
        spike_out_source422 = spike_out_source_array[422];
    end
    always @(spike_out_source_array[423]) begin 
        spike_out_source423 = spike_out_source_array[423];
    end
    always @(spike_out_source_array[424]) begin 
        spike_out_source424 = spike_out_source_array[424];
    end
    always @(spike_out_source_array[425]) begin 
        spike_out_source425 = spike_out_source_array[425];
    end
    always @(spike_out_source_array[426]) begin 
        spike_out_source426 = spike_out_source_array[426];
    end
    always @(spike_out_source_array[427]) begin 
        spike_out_source427 = spike_out_source_array[427];
    end
    always @(spike_out_source_array[428]) begin 
        spike_out_source428 = spike_out_source_array[428];
    end
    always @(spike_out_source_array[429]) begin 
        spike_out_source429 = spike_out_source_array[429];
    end
    always @(spike_out_source_array[430]) begin 
        spike_out_source430 = spike_out_source_array[430];
    end
    always @(spike_out_source_array[431]) begin 
        spike_out_source431 = spike_out_source_array[431];
    end
    always @(spike_out_source_array[432]) begin 
        spike_out_source432 = spike_out_source_array[432];
    end
    always @(spike_out_source_array[433]) begin 
        spike_out_source433 = spike_out_source_array[433];
    end
    always @(spike_out_source_array[434]) begin 
        spike_out_source434 = spike_out_source_array[434];
    end
    always @(spike_out_source_array[435]) begin 
        spike_out_source435 = spike_out_source_array[435];
    end
    always @(spike_out_source_array[436]) begin 
        spike_out_source436 = spike_out_source_array[436];
    end
    always @(spike_out_source_array[437]) begin 
        spike_out_source437 = spike_out_source_array[437];
    end
    always @(spike_out_source_array[438]) begin 
        spike_out_source438 = spike_out_source_array[438];
    end
    always @(spike_out_source_array[439]) begin 
        spike_out_source439 = spike_out_source_array[439];
    end
    always @(spike_out_source_array[440]) begin 
        spike_out_source440 = spike_out_source_array[440];
    end
    always @(spike_out_source_array[441]) begin 
        spike_out_source441 = spike_out_source_array[441];
    end
    always @(spike_out_source_array[442]) begin 
        spike_out_source442 = spike_out_source_array[442];
    end
    always @(spike_out_source_array[443]) begin 
        spike_out_source443 = spike_out_source_array[443];
    end
    always @(spike_out_source_array[444]) begin 
        spike_out_source444 = spike_out_source_array[444];
    end
    always @(spike_out_source_array[445]) begin 
        spike_out_source445 = spike_out_source_array[445];
    end
    always @(spike_out_source_array[446]) begin 
        spike_out_source446 = spike_out_source_array[446];
    end
    always @(spike_out_source_array[447]) begin 
        spike_out_source447 = spike_out_source_array[447];
    end
    always @(spike_out_source_array[448]) begin 
        spike_out_source448 = spike_out_source_array[448];
    end
    always @(spike_out_source_array[449]) begin 
        spike_out_source449 = spike_out_source_array[449];
    end
    always @(spike_out_source_array[450]) begin 
        spike_out_source450 = spike_out_source_array[450];
    end
    always @(spike_out_source_array[451]) begin 
        spike_out_source451 = spike_out_source_array[451];
    end
    always @(spike_out_source_array[452]) begin 
        spike_out_source452 = spike_out_source_array[452];
    end
    always @(spike_out_source_array[453]) begin 
        spike_out_source453 = spike_out_source_array[453];
    end
    always @(spike_out_source_array[454]) begin 
        spike_out_source454 = spike_out_source_array[454];
    end
    always @(spike_out_source_array[455]) begin 
        spike_out_source455 = spike_out_source_array[455];
    end
    always @(spike_out_source_array[456]) begin 
        spike_out_source456 = spike_out_source_array[456];
    end
    always @(spike_out_source_array[457]) begin 
        spike_out_source457 = spike_out_source_array[457];
    end
    always @(spike_out_source_array[458]) begin 
        spike_out_source458 = spike_out_source_array[458];
    end
    always @(spike_out_source_array[459]) begin 
        spike_out_source459 = spike_out_source_array[459];
    end
    always @(spike_out_source_array[460]) begin 
        spike_out_source460 = spike_out_source_array[460];
    end
    always @(spike_out_source_array[461]) begin 
        spike_out_source461 = spike_out_source_array[461];
    end
    always @(spike_out_source_array[462]) begin 
        spike_out_source462 = spike_out_source_array[462];
    end
    always @(spike_out_source_array[463]) begin 
        spike_out_source463 = spike_out_source_array[463];
    end
    always @(spike_out_source_array[464]) begin 
        spike_out_source464 = spike_out_source_array[464];
    end
    always @(spike_out_source_array[465]) begin 
        spike_out_source465 = spike_out_source_array[465];
    end
    always @(spike_out_source_array[466]) begin 
        spike_out_source466 = spike_out_source_array[466];
    end
    always @(spike_out_source_array[467]) begin 
        spike_out_source467 = spike_out_source_array[467];
    end
    always @(spike_out_source_array[468]) begin 
        spike_out_source468 = spike_out_source_array[468];
    end
    always @(spike_out_source_array[469]) begin 
        spike_out_source469 = spike_out_source_array[469];
    end
    always @(spike_out_source_array[470]) begin 
        spike_out_source470 = spike_out_source_array[470];
    end
    always @(spike_out_source_array[471]) begin 
        spike_out_source471 = spike_out_source_array[471];
    end
    always @(spike_out_source_array[472]) begin 
        spike_out_source472 = spike_out_source_array[472];
    end
    always @(spike_out_source_array[473]) begin 
        spike_out_source473 = spike_out_source_array[473];
    end
    always @(spike_out_source_array[474]) begin 
        spike_out_source474 = spike_out_source_array[474];
    end
    always @(spike_out_source_array[475]) begin 
        spike_out_source475 = spike_out_source_array[475];
    end
    always @(spike_out_source_array[476]) begin 
        spike_out_source476 = spike_out_source_array[476];
    end
    always @(spike_out_source_array[477]) begin 
        spike_out_source477 = spike_out_source_array[477];
    end
    always @(spike_out_source_array[478]) begin 
        spike_out_source478 = spike_out_source_array[478];
    end
    always @(spike_out_source_array[479]) begin 
        spike_out_source479 = spike_out_source_array[479];
    end
    always @(spike_out_source_array[480]) begin 
        spike_out_source480 = spike_out_source_array[480];
    end
    always @(spike_out_source_array[481]) begin 
        spike_out_source481 = spike_out_source_array[481];
    end
    always @(spike_out_source_array[482]) begin 
        spike_out_source482 = spike_out_source_array[482];
    end
    always @(spike_out_source_array[483]) begin 
        spike_out_source483 = spike_out_source_array[483];
    end
    always @(spike_out_source_array[484]) begin 
        spike_out_source484 = spike_out_source_array[484];
    end
    always @(spike_out_source_array[485]) begin 
        spike_out_source485 = spike_out_source_array[485];
    end
    always @(spike_out_source_array[486]) begin 
        spike_out_source486 = spike_out_source_array[486];
    end
    always @(spike_out_source_array[487]) begin 
        spike_out_source487 = spike_out_source_array[487];
    end
    always @(spike_out_source_array[488]) begin 
        spike_out_source488 = spike_out_source_array[488];
    end
    always @(spike_out_source_array[489]) begin 
        spike_out_source489 = spike_out_source_array[489];
    end
    always @(spike_out_source_array[490]) begin 
        spike_out_source490 = spike_out_source_array[490];
    end
    always @(spike_out_source_array[491]) begin 
        spike_out_source491 = spike_out_source_array[491];
    end
    always @(spike_out_source_array[492]) begin 
        spike_out_source492 = spike_out_source_array[492];
    end
    always @(spike_out_source_array[493]) begin 
        spike_out_source493 = spike_out_source_array[493];
    end
    always @(spike_out_source_array[494]) begin 
        spike_out_source494 = spike_out_source_array[494];
    end
    always @(spike_out_source_array[495]) begin 
        spike_out_source495 = spike_out_source_array[495];
    end
    always @(spike_out_source_array[496]) begin 
        spike_out_source496 = spike_out_source_array[496];
    end
    always @(spike_out_source_array[497]) begin 
        spike_out_source497 = spike_out_source_array[497];
    end
    always @(spike_out_source_array[498]) begin 
        spike_out_source498 = spike_out_source_array[498];
    end
    always @(spike_out_source_array[499]) begin 
        spike_out_source499 = spike_out_source_array[499];
    end
    always @(spike_out_source_array[500]) begin 
        spike_out_source500 = spike_out_source_array[500];
    end
    always @(spike_out_source_array[501]) begin 
        spike_out_source501 = spike_out_source_array[501];
    end
    always @(spike_out_source_array[502]) begin 
        spike_out_source502 = spike_out_source_array[502];
    end
    always @(spike_out_source_array[503]) begin 
        spike_out_source503 = spike_out_source_array[503];
    end
    always @(spike_out_source_array[504]) begin 
        spike_out_source504 = spike_out_source_array[504];
    end
    always @(spike_out_source_array[505]) begin 
        spike_out_source505 = spike_out_source_array[505];
    end
    always @(spike_out_source_array[506]) begin 
        spike_out_source506 = spike_out_source_array[506];
    end
    always @(spike_out_source_array[507]) begin 
        spike_out_source507 = spike_out_source_array[507];
    end
    always @(spike_out_source_array[508]) begin 
        spike_out_source508 = spike_out_source_array[508];
    end
    always @(spike_out_source_array[509]) begin 
        spike_out_source509 = spike_out_source_array[509];
    end
    always @(spike_out_source_array[510]) begin 
        spike_out_source510 = spike_out_source_array[510];
    end
    always @(spike_out_source_array[511]) begin 
        spike_out_source511 = spike_out_source_array[511];
    end
    always @(spike_out_source_array[512]) begin 
        spike_out_source512 = spike_out_source_array[512];
    end
    always @(spike_out_source_array[513]) begin 
        spike_out_source513 = spike_out_source_array[513];
    end
    always @(spike_out_source_array[514]) begin 
        spike_out_source514 = spike_out_source_array[514];
    end
    always @(spike_out_source_array[515]) begin 
        spike_out_source515 = spike_out_source_array[515];
    end
    always @(spike_out_source_array[516]) begin 
        spike_out_source516 = spike_out_source_array[516];
    end
    always @(spike_out_source_array[517]) begin 
        spike_out_source517 = spike_out_source_array[517];
    end
    always @(spike_out_source_array[518]) begin 
        spike_out_source518 = spike_out_source_array[518];
    end
    always @(spike_out_source_array[519]) begin 
        spike_out_source519 = spike_out_source_array[519];
    end
    always @(spike_out_source_array[520]) begin 
        spike_out_source520 = spike_out_source_array[520];
    end
    always @(spike_out_source_array[521]) begin 
        spike_out_source521 = spike_out_source_array[521];
    end
    always @(spike_out_source_array[522]) begin 
        spike_out_source522 = spike_out_source_array[522];
    end
    always @(spike_out_source_array[523]) begin 
        spike_out_source523 = spike_out_source_array[523];
    end
    always @(spike_out_source_array[524]) begin 
        spike_out_source524 = spike_out_source_array[524];
    end
    always @(spike_out_source_array[525]) begin 
        spike_out_source525 = spike_out_source_array[525];
    end
    always @(spike_out_source_array[526]) begin 
        spike_out_source526 = spike_out_source_array[526];
    end
    always @(spike_out_source_array[527]) begin 
        spike_out_source527 = spike_out_source_array[527];
    end
    always @(spike_out_source_array[528]) begin 
        spike_out_source528 = spike_out_source_array[528];
    end
    always @(spike_out_source_array[529]) begin 
        spike_out_source529 = spike_out_source_array[529];
    end
    always @(spike_out_source_array[530]) begin 
        spike_out_source530 = spike_out_source_array[530];
    end
    always @(spike_out_source_array[531]) begin 
        spike_out_source531 = spike_out_source_array[531];
    end
    always @(spike_out_source_array[532]) begin 
        spike_out_source532 = spike_out_source_array[532];
    end
    always @(spike_out_source_array[533]) begin 
        spike_out_source533 = spike_out_source_array[533];
    end
    always @(spike_out_source_array[534]) begin 
        spike_out_source534 = spike_out_source_array[534];
    end
    always @(spike_out_source_array[535]) begin 
        spike_out_source535 = spike_out_source_array[535];
    end
    always @(spike_out_source_array[536]) begin 
        spike_out_source536 = spike_out_source_array[536];
    end
    always @(spike_out_source_array[537]) begin 
        spike_out_source537 = spike_out_source_array[537];
    end
    always @(spike_out_source_array[538]) begin 
        spike_out_source538 = spike_out_source_array[538];
    end
    always @(spike_out_source_array[539]) begin 
        spike_out_source539 = spike_out_source_array[539];
    end
    always @(spike_out_source_array[540]) begin 
        spike_out_source540 = spike_out_source_array[540];
    end
    always @(spike_out_source_array[541]) begin 
        spike_out_source541 = spike_out_source_array[541];
    end
    always @(spike_out_source_array[542]) begin 
        spike_out_source542 = spike_out_source_array[542];
    end
    always @(spike_out_source_array[543]) begin 
        spike_out_source543 = spike_out_source_array[543];
    end
    always @(spike_out_source_array[544]) begin 
        spike_out_source544 = spike_out_source_array[544];
    end
    always @(spike_out_source_array[545]) begin 
        spike_out_source545 = spike_out_source_array[545];
    end
    always @(spike_out_source_array[546]) begin 
        spike_out_source546 = spike_out_source_array[546];
    end
    always @(spike_out_source_array[547]) begin 
        spike_out_source547 = spike_out_source_array[547];
    end
    always @(spike_out_source_array[548]) begin 
        spike_out_source548 = spike_out_source_array[548];
    end
    always @(spike_out_source_array[549]) begin 
        spike_out_source549 = spike_out_source_array[549];
    end
    always @(spike_out_source_array[550]) begin 
        spike_out_source550 = spike_out_source_array[550];
    end
    always @(spike_out_source_array[551]) begin 
        spike_out_source551 = spike_out_source_array[551];
    end
    always @(spike_out_source_array[552]) begin 
        spike_out_source552 = spike_out_source_array[552];
    end
    always @(spike_out_source_array[553]) begin 
        spike_out_source553 = spike_out_source_array[553];
    end
    always @(spike_out_source_array[554]) begin 
        spike_out_source554 = spike_out_source_array[554];
    end
    always @(spike_out_source_array[555]) begin 
        spike_out_source555 = spike_out_source_array[555];
    end
    always @(spike_out_source_array[556]) begin 
        spike_out_source556 = spike_out_source_array[556];
    end
    always @(spike_out_source_array[557]) begin 
        spike_out_source557 = spike_out_source_array[557];
    end
    always @(spike_out_source_array[558]) begin 
        spike_out_source558 = spike_out_source_array[558];
    end
    always @(spike_out_source_array[559]) begin 
        spike_out_source559 = spike_out_source_array[559];
    end
    always @(spike_out_source_array[560]) begin 
        spike_out_source560 = spike_out_source_array[560];
    end
    always @(spike_out_source_array[561]) begin 
        spike_out_source561 = spike_out_source_array[561];
    end
    always @(spike_out_source_array[562]) begin 
        spike_out_source562 = spike_out_source_array[562];
    end
    always @(spike_out_source_array[563]) begin 
        spike_out_source563 = spike_out_source_array[563];
    end
    always @(spike_out_source_array[564]) begin 
        spike_out_source564 = spike_out_source_array[564];
    end
    always @(spike_out_source_array[565]) begin 
        spike_out_source565 = spike_out_source_array[565];
    end
    always @(spike_out_source_array[566]) begin 
        spike_out_source566 = spike_out_source_array[566];
    end
    always @(spike_out_source_array[567]) begin 
        spike_out_source567 = spike_out_source_array[567];
    end
    always @(spike_out_source_array[568]) begin 
        spike_out_source568 = spike_out_source_array[568];
    end
    always @(spike_out_source_array[569]) begin 
        spike_out_source569 = spike_out_source_array[569];
    end
    always @(spike_out_source_array[570]) begin 
        spike_out_source570 = spike_out_source_array[570];
    end
    always @(spike_out_source_array[571]) begin 
        spike_out_source571 = spike_out_source_array[571];
    end
    always @(spike_out_source_array[572]) begin 
        spike_out_source572 = spike_out_source_array[572];
    end
    always @(spike_out_source_array[573]) begin 
        spike_out_source573 = spike_out_source_array[573];
    end
    always @(spike_out_source_array[574]) begin 
        spike_out_source574 = spike_out_source_array[574];
    end
    always @(spike_out_source_array[575]) begin 
        spike_out_source575 = spike_out_source_array[575];
    end
    always @(spike_out_source_array[576]) begin 
        spike_out_source576 = spike_out_source_array[576];
    end
    always @(spike_out_source_array[577]) begin 
        spike_out_source577 = spike_out_source_array[577];
    end
    always @(spike_out_source_array[578]) begin 
        spike_out_source578 = spike_out_source_array[578];
    end
    always @(spike_out_source_array[579]) begin 
        spike_out_source579 = spike_out_source_array[579];
    end
    always @(spike_out_source_array[580]) begin 
        spike_out_source580 = spike_out_source_array[580];
    end
    always @(spike_out_source_array[581]) begin 
        spike_out_source581 = spike_out_source_array[581];
    end
    always @(spike_out_source_array[582]) begin 
        spike_out_source582 = spike_out_source_array[582];
    end
    always @(spike_out_source_array[583]) begin 
        spike_out_source583 = spike_out_source_array[583];
    end
    always @(spike_out_source_array[584]) begin 
        spike_out_source584 = spike_out_source_array[584];
    end
    always @(spike_out_source_array[585]) begin 
        spike_out_source585 = spike_out_source_array[585];
    end
    always @(spike_out_source_array[586]) begin 
        spike_out_source586 = spike_out_source_array[586];
    end
    always @(spike_out_source_array[587]) begin 
        spike_out_source587 = spike_out_source_array[587];
    end
    always @(spike_out_source_array[588]) begin 
        spike_out_source588 = spike_out_source_array[588];
    end
    always @(spike_out_source_array[589]) begin 
        spike_out_source589 = spike_out_source_array[589];
    end
    always @(spike_out_source_array[590]) begin 
        spike_out_source590 = spike_out_source_array[590];
    end
    always @(spike_out_source_array[591]) begin 
        spike_out_source591 = spike_out_source_array[591];
    end
    always @(spike_out_source_array[592]) begin 
        spike_out_source592 = spike_out_source_array[592];
    end
    always @(spike_out_source_array[593]) begin 
        spike_out_source593 = spike_out_source_array[593];
    end
    always @(spike_out_source_array[594]) begin 
        spike_out_source594 = spike_out_source_array[594];
    end
    always @(spike_out_source_array[595]) begin 
        spike_out_source595 = spike_out_source_array[595];
    end
    always @(spike_out_source_array[596]) begin 
        spike_out_source596 = spike_out_source_array[596];
    end
    always @(spike_out_source_array[597]) begin 
        spike_out_source597 = spike_out_source_array[597];
    end
    always @(spike_out_source_array[598]) begin 
        spike_out_source598 = spike_out_source_array[598];
    end
    always @(spike_out_source_array[599]) begin 
        spike_out_source599 = spike_out_source_array[599];
    end
    always @(spike_out_source_array[600]) begin 
        spike_out_source600 = spike_out_source_array[600];
    end
    always @(spike_out_source_array[601]) begin 
        spike_out_source601 = spike_out_source_array[601];
    end
    always @(spike_out_source_array[602]) begin 
        spike_out_source602 = spike_out_source_array[602];
    end
    always @(spike_out_source_array[603]) begin 
        spike_out_source603 = spike_out_source_array[603];
    end
    always @(spike_out_source_array[604]) begin 
        spike_out_source604 = spike_out_source_array[604];
    end
    always @(spike_out_source_array[605]) begin 
        spike_out_source605 = spike_out_source_array[605];
    end
    always @(spike_out_source_array[606]) begin 
        spike_out_source606 = spike_out_source_array[606];
    end
    always @(spike_out_source_array[607]) begin 
        spike_out_source607 = spike_out_source_array[607];
    end
    always @(spike_out_source_array[608]) begin 
        spike_out_source608 = spike_out_source_array[608];
    end
    always @(spike_out_source_array[609]) begin 
        spike_out_source609 = spike_out_source_array[609];
    end
    always @(spike_out_source_array[610]) begin 
        spike_out_source610 = spike_out_source_array[610];
    end
    always @(spike_out_source_array[611]) begin 
        spike_out_source611 = spike_out_source_array[611];
    end
    always @(spike_out_source_array[612]) begin 
        spike_out_source612 = spike_out_source_array[612];
    end
    always @(spike_out_source_array[613]) begin 
        spike_out_source613 = spike_out_source_array[613];
    end
    always @(spike_out_source_array[614]) begin 
        spike_out_source614 = spike_out_source_array[614];
    end
    always @(spike_out_source_array[615]) begin 
        spike_out_source615 = spike_out_source_array[615];
    end
    always @(spike_out_source_array[616]) begin 
        spike_out_source616 = spike_out_source_array[616];
    end
    always @(spike_out_source_array[617]) begin 
        spike_out_source617 = spike_out_source_array[617];
    end
    always @(spike_out_source_array[618]) begin 
        spike_out_source618 = spike_out_source_array[618];
    end
    always @(spike_out_source_array[619]) begin 
        spike_out_source619 = spike_out_source_array[619];
    end
    always @(spike_out_source_array[620]) begin 
        spike_out_source620 = spike_out_source_array[620];
    end
    always @(spike_out_source_array[621]) begin 
        spike_out_source621 = spike_out_source_array[621];
    end
    always @(spike_out_source_array[622]) begin 
        spike_out_source622 = spike_out_source_array[622];
    end
    always @(spike_out_source_array[623]) begin 
        spike_out_source623 = spike_out_source_array[623];
    end
    always @(spike_out_source_array[624]) begin 
        spike_out_source624 = spike_out_source_array[624];
    end
    always @(spike_out_source_array[625]) begin 
        spike_out_source625 = spike_out_source_array[625];
    end
    always @(spike_out_source_array[626]) begin 
        spike_out_source626 = spike_out_source_array[626];
    end
    always @(spike_out_source_array[627]) begin 
        spike_out_source627 = spike_out_source_array[627];
    end
    always @(spike_out_source_array[628]) begin 
        spike_out_source628 = spike_out_source_array[628];
    end
    always @(spike_out_source_array[629]) begin 
        spike_out_source629 = spike_out_source_array[629];
    end
    always @(spike_out_source_array[630]) begin 
        spike_out_source630 = spike_out_source_array[630];
    end
    always @(spike_out_source_array[631]) begin 
        spike_out_source631 = spike_out_source_array[631];
    end
    always @(spike_out_source_array[632]) begin 
        spike_out_source632 = spike_out_source_array[632];
    end
    always @(spike_out_source_array[633]) begin 
        spike_out_source633 = spike_out_source_array[633];
    end
    always @(spike_out_source_array[634]) begin 
        spike_out_source634 = spike_out_source_array[634];
    end
    always @(spike_out_source_array[635]) begin 
        spike_out_source635 = spike_out_source_array[635];
    end
    always @(spike_out_source_array[636]) begin 
        spike_out_source636 = spike_out_source_array[636];
    end
    always @(spike_out_source_array[637]) begin 
        spike_out_source637 = spike_out_source_array[637];
    end
    always @(spike_out_source_array[638]) begin 
        spike_out_source638 = spike_out_source_array[638];
    end
    always @(spike_out_source_array[639]) begin 
        spike_out_source639 = spike_out_source_array[639];
    end
    always @(spike_out_source_array[640]) begin 
        spike_out_source640 = spike_out_source_array[640];
    end
    always @(spike_out_source_array[641]) begin 
        spike_out_source641 = spike_out_source_array[641];
    end
    always @(spike_out_source_array[642]) begin 
        spike_out_source642 = spike_out_source_array[642];
    end
    always @(spike_out_source_array[643]) begin 
        spike_out_source643 = spike_out_source_array[643];
    end
    always @(spike_out_source_array[644]) begin 
        spike_out_source644 = spike_out_source_array[644];
    end
    always @(spike_out_source_array[645]) begin 
        spike_out_source645 = spike_out_source_array[645];
    end
    always @(spike_out_source_array[646]) begin 
        spike_out_source646 = spike_out_source_array[646];
    end
    always @(spike_out_source_array[647]) begin 
        spike_out_source647 = spike_out_source_array[647];
    end
    always @(spike_out_source_array[648]) begin 
        spike_out_source648 = spike_out_source_array[648];
    end
    always @(spike_out_source_array[649]) begin 
        spike_out_source649 = spike_out_source_array[649];
    end
    always @(spike_out_source_array[650]) begin 
        spike_out_source650 = spike_out_source_array[650];
    end
    always @(spike_out_source_array[651]) begin 
        spike_out_source651 = spike_out_source_array[651];
    end
    always @(spike_out_source_array[652]) begin 
        spike_out_source652 = spike_out_source_array[652];
    end
    always @(spike_out_source_array[653]) begin 
        spike_out_source653 = spike_out_source_array[653];
    end
    always @(spike_out_source_array[654]) begin 
        spike_out_source654 = spike_out_source_array[654];
    end
    always @(spike_out_source_array[655]) begin 
        spike_out_source655 = spike_out_source_array[655];
    end
    always @(spike_out_source_array[656]) begin 
        spike_out_source656 = spike_out_source_array[656];
    end
    always @(spike_out_source_array[657]) begin 
        spike_out_source657 = spike_out_source_array[657];
    end
    always @(spike_out_source_array[658]) begin 
        spike_out_source658 = spike_out_source_array[658];
    end
    always @(spike_out_source_array[659]) begin 
        spike_out_source659 = spike_out_source_array[659];
    end
    always @(spike_out_source_array[660]) begin 
        spike_out_source660 = spike_out_source_array[660];
    end
    always @(spike_out_source_array[661]) begin 
        spike_out_source661 = spike_out_source_array[661];
    end
    always @(spike_out_source_array[662]) begin 
        spike_out_source662 = spike_out_source_array[662];
    end
    always @(spike_out_source_array[663]) begin 
        spike_out_source663 = spike_out_source_array[663];
    end
    always @(spike_out_source_array[664]) begin 
        spike_out_source664 = spike_out_source_array[664];
    end
    always @(spike_out_source_array[665]) begin 
        spike_out_source665 = spike_out_source_array[665];
    end
    always @(spike_out_source_array[666]) begin 
        spike_out_source666 = spike_out_source_array[666];
    end
    always @(spike_out_source_array[667]) begin 
        spike_out_source667 = spike_out_source_array[667];
    end
    always @(spike_out_source_array[668]) begin 
        spike_out_source668 = spike_out_source_array[668];
    end
    always @(spike_out_source_array[669]) begin 
        spike_out_source669 = spike_out_source_array[669];
    end
    always @(spike_out_source_array[670]) begin 
        spike_out_source670 = spike_out_source_array[670];
    end
    always @(spike_out_source_array[671]) begin 
        spike_out_source671 = spike_out_source_array[671];
    end
    always @(spike_out_source_array[672]) begin 
        spike_out_source672 = spike_out_source_array[672];
    end
    always @(spike_out_source_array[673]) begin 
        spike_out_source673 = spike_out_source_array[673];
    end
    always @(spike_out_source_array[674]) begin 
        spike_out_source674 = spike_out_source_array[674];
    end
    always @(spike_out_source_array[675]) begin 
        spike_out_source675 = spike_out_source_array[675];
    end
    always @(spike_out_source_array[676]) begin 
        spike_out_source676 = spike_out_source_array[676];
    end
    always @(spike_out_source_array[677]) begin 
        spike_out_source677 = spike_out_source_array[677];
    end
    always @(spike_out_source_array[678]) begin 
        spike_out_source678 = spike_out_source_array[678];
    end
    always @(spike_out_source_array[679]) begin 
        spike_out_source679 = spike_out_source_array[679];
    end
    always @(spike_out_source_array[680]) begin 
        spike_out_source680 = spike_out_source_array[680];
    end
    always @(spike_out_source_array[681]) begin 
        spike_out_source681 = spike_out_source_array[681];
    end
    always @(spike_out_source_array[682]) begin 
        spike_out_source682 = spike_out_source_array[682];
    end
    always @(spike_out_source_array[683]) begin 
        spike_out_source683 = spike_out_source_array[683];
    end
    always @(spike_out_source_array[684]) begin 
        spike_out_source684 = spike_out_source_array[684];
    end
    always @(spike_out_source_array[685]) begin 
        spike_out_source685 = spike_out_source_array[685];
    end
    always @(spike_out_source_array[686]) begin 
        spike_out_source686 = spike_out_source_array[686];
    end
    always @(spike_out_source_array[687]) begin 
        spike_out_source687 = spike_out_source_array[687];
    end
    always @(spike_out_source_array[688]) begin 
        spike_out_source688 = spike_out_source_array[688];
    end
    always @(spike_out_source_array[689]) begin 
        spike_out_source689 = spike_out_source_array[689];
    end
    always @(spike_out_source_array[690]) begin 
        spike_out_source690 = spike_out_source_array[690];
    end
    always @(spike_out_source_array[691]) begin 
        spike_out_source691 = spike_out_source_array[691];
    end
    always @(spike_out_source_array[692]) begin 
        spike_out_source692 = spike_out_source_array[692];
    end
    always @(spike_out_source_array[693]) begin 
        spike_out_source693 = spike_out_source_array[693];
    end
    always @(spike_out_source_array[694]) begin 
        spike_out_source694 = spike_out_source_array[694];
    end
    always @(spike_out_source_array[695]) begin 
        spike_out_source695 = spike_out_source_array[695];
    end
    always @(spike_out_source_array[696]) begin 
        spike_out_source696 = spike_out_source_array[696];
    end
    always @(spike_out_source_array[697]) begin 
        spike_out_source697 = spike_out_source_array[697];
    end
    always @(spike_out_source_array[698]) begin 
        spike_out_source698 = spike_out_source_array[698];
    end
    always @(spike_out_source_array[699]) begin 
        spike_out_source699 = spike_out_source_array[699];
    end
    always @(spike_out_source_array[700]) begin 
        spike_out_source700 = spike_out_source_array[700];
    end
    always @(spike_out_source_array[701]) begin 
        spike_out_source701 = spike_out_source_array[701];
    end
    always @(spike_out_source_array[702]) begin 
        spike_out_source702 = spike_out_source_array[702];
    end
    always @(spike_out_source_array[703]) begin 
        spike_out_source703 = spike_out_source_array[703];
    end
    always @(spike_out_source_array[704]) begin 
        spike_out_source704 = spike_out_source_array[704];
    end
    always @(spike_out_source_array[705]) begin 
        spike_out_source705 = spike_out_source_array[705];
    end
    always @(spike_out_source_array[706]) begin 
        spike_out_source706 = spike_out_source_array[706];
    end
    always @(spike_out_source_array[707]) begin 
        spike_out_source707 = spike_out_source_array[707];
    end
    always @(spike_out_source_array[708]) begin 
        spike_out_source708 = spike_out_source_array[708];
    end
    always @(spike_out_source_array[709]) begin 
        spike_out_source709 = spike_out_source_array[709];
    end
    always @(spike_out_source_array[710]) begin 
        spike_out_source710 = spike_out_source_array[710];
    end
    always @(spike_out_source_array[711]) begin 
        spike_out_source711 = spike_out_source_array[711];
    end
    always @(spike_out_source_array[712]) begin 
        spike_out_source712 = spike_out_source_array[712];
    end
    always @(spike_out_source_array[713]) begin 
        spike_out_source713 = spike_out_source_array[713];
    end
    always @(spike_out_source_array[714]) begin 
        spike_out_source714 = spike_out_source_array[714];
    end
    always @(spike_out_source_array[715]) begin 
        spike_out_source715 = spike_out_source_array[715];
    end
    always @(spike_out_source_array[716]) begin 
        spike_out_source716 = spike_out_source_array[716];
    end
    always @(spike_out_source_array[717]) begin 
        spike_out_source717 = spike_out_source_array[717];
    end
    always @(spike_out_source_array[718]) begin 
        spike_out_source718 = spike_out_source_array[718];
    end
    always @(spike_out_source_array[719]) begin 
        spike_out_source719 = spike_out_source_array[719];
    end
    always @(spike_out_source_array[720]) begin 
        spike_out_source720 = spike_out_source_array[720];
    end
    always @(spike_out_source_array[721]) begin 
        spike_out_source721 = spike_out_source_array[721];
    end
    always @(spike_out_source_array[722]) begin 
        spike_out_source722 = spike_out_source_array[722];
    end
    always @(spike_out_source_array[723]) begin 
        spike_out_source723 = spike_out_source_array[723];
    end
    always @(spike_out_source_array[724]) begin 
        spike_out_source724 = spike_out_source_array[724];
    end
    always @(spike_out_source_array[725]) begin 
        spike_out_source725 = spike_out_source_array[725];
    end
    always @(spike_out_source_array[726]) begin 
        spike_out_source726 = spike_out_source_array[726];
    end
    always @(spike_out_source_array[727]) begin 
        spike_out_source727 = spike_out_source_array[727];
    end
    always @(spike_out_source_array[728]) begin 
        spike_out_source728 = spike_out_source_array[728];
    end
    always @(spike_out_source_array[729]) begin 
        spike_out_source729 = spike_out_source_array[729];
    end
    always @(spike_out_source_array[730]) begin 
        spike_out_source730 = spike_out_source_array[730];
    end
    always @(spike_out_source_array[731]) begin 
        spike_out_source731 = spike_out_source_array[731];
    end
    always @(spike_out_source_array[732]) begin 
        spike_out_source732 = spike_out_source_array[732];
    end
    always @(spike_out_source_array[733]) begin 
        spike_out_source733 = spike_out_source_array[733];
    end
    always @(spike_out_source_array[734]) begin 
        spike_out_source734 = spike_out_source_array[734];
    end
    always @(spike_out_source_array[735]) begin 
        spike_out_source735 = spike_out_source_array[735];
    end
    always @(spike_out_source_array[736]) begin 
        spike_out_source736 = spike_out_source_array[736];
    end
    always @(spike_out_source_array[737]) begin 
        spike_out_source737 = spike_out_source_array[737];
    end
    always @(spike_out_source_array[738]) begin 
        spike_out_source738 = spike_out_source_array[738];
    end
    always @(spike_out_source_array[739]) begin 
        spike_out_source739 = spike_out_source_array[739];
    end
    always @(spike_out_source_array[740]) begin 
        spike_out_source740 = spike_out_source_array[740];
    end
    always @(spike_out_source_array[741]) begin 
        spike_out_source741 = spike_out_source_array[741];
    end
    always @(spike_out_source_array[742]) begin 
        spike_out_source742 = spike_out_source_array[742];
    end
    always @(spike_out_source_array[743]) begin 
        spike_out_source743 = spike_out_source_array[743];
    end
    always @(spike_out_source_array[744]) begin 
        spike_out_source744 = spike_out_source_array[744];
    end
    always @(spike_out_source_array[745]) begin 
        spike_out_source745 = spike_out_source_array[745];
    end
    always @(spike_out_source_array[746]) begin 
        spike_out_source746 = spike_out_source_array[746];
    end
    always @(spike_out_source_array[747]) begin 
        spike_out_source747 = spike_out_source_array[747];
    end
    always @(spike_out_source_array[748]) begin 
        spike_out_source748 = spike_out_source_array[748];
    end
    always @(spike_out_source_array[749]) begin 
        spike_out_source749 = spike_out_source_array[749];
    end
    always @(spike_out_source_array[750]) begin 
        spike_out_source750 = spike_out_source_array[750];
    end
    always @(spike_out_source_array[751]) begin 
        spike_out_source751 = spike_out_source_array[751];
    end
    always @(spike_out_source_array[752]) begin 
        spike_out_source752 = spike_out_source_array[752];
    end
    always @(spike_out_source_array[753]) begin 
        spike_out_source753 = spike_out_source_array[753];
    end
    always @(spike_out_source_array[754]) begin 
        spike_out_source754 = spike_out_source_array[754];
    end
    always @(spike_out_source_array[755]) begin 
        spike_out_source755 = spike_out_source_array[755];
    end
    always @(spike_out_source_array[756]) begin 
        spike_out_source756 = spike_out_source_array[756];
    end
    always @(spike_out_source_array[757]) begin 
        spike_out_source757 = spike_out_source_array[757];
    end
    always @(spike_out_source_array[758]) begin 
        spike_out_source758 = spike_out_source_array[758];
    end
    always @(spike_out_source_array[759]) begin 
        spike_out_source759 = spike_out_source_array[759];
    end
    always @(spike_out_source_array[760]) begin 
        spike_out_source760 = spike_out_source_array[760];
    end
    always @(spike_out_source_array[761]) begin 
        spike_out_source761 = spike_out_source_array[761];
    end
    always @(spike_out_source_array[762]) begin 
        spike_out_source762 = spike_out_source_array[762];
    end
    always @(spike_out_source_array[763]) begin 
        spike_out_source763 = spike_out_source_array[763];
    end
    always @(spike_out_source_array[764]) begin 
        spike_out_source764 = spike_out_source_array[764];
    end
    always @(spike_out_source_array[765]) begin 
        spike_out_source765 = spike_out_source_array[765];
    end
    always @(spike_out_source_array[766]) begin 
        spike_out_source766 = spike_out_source_array[766];
    end
    always @(spike_out_source_array[767]) begin 
        spike_out_source767 = spike_out_source_array[767];
    end
    always @(spike_out_source_array[768]) begin 
        spike_out_source768 = spike_out_source_array[768];
    end
    always @(spike_out_source_array[769]) begin 
        spike_out_source769 = spike_out_source_array[769];
    end
    always @(spike_out_source_array[770]) begin 
        spike_out_source770 = spike_out_source_array[770];
    end
    always @(spike_out_source_array[771]) begin 
        spike_out_source771 = spike_out_source_array[771];
    end
    always @(spike_out_source_array[772]) begin 
        spike_out_source772 = spike_out_source_array[772];
    end
    always @(spike_out_source_array[773]) begin 
        spike_out_source773 = spike_out_source_array[773];
    end
    always @(spike_out_source_array[774]) begin 
        spike_out_source774 = spike_out_source_array[774];
    end
    always @(spike_out_source_array[775]) begin 
        spike_out_source775 = spike_out_source_array[775];
    end
    always @(spike_out_source_array[776]) begin 
        spike_out_source776 = spike_out_source_array[776];
    end
    always @(spike_out_source_array[777]) begin 
        spike_out_source777 = spike_out_source_array[777];
    end
    always @(spike_out_source_array[778]) begin 
        spike_out_source778 = spike_out_source_array[778];
    end
    always @(spike_out_source_array[779]) begin 
        spike_out_source779 = spike_out_source_array[779];
    end
    always @(spike_out_source_array[780]) begin 
        spike_out_source780 = spike_out_source_array[780];
    end
    always @(spike_out_source_array[781]) begin 
        spike_out_source781 = spike_out_source_array[781];
    end
    always @(spike_out_source_array[782]) begin 
        spike_out_source782 = spike_out_source_array[782];
    end
    always @(spike_out_source_array[783]) begin 
        spike_out_source783 = spike_out_source_array[783];
    end
    always @(spike_out_source_array[784]) begin 
        spike_out_source784 = spike_out_source_array[784];
    end
    always @(spike_out_source_array[785]) begin 
        spike_out_source785 = spike_out_source_array[785];
    end
    always @(spike_out_source_array[786]) begin 
        spike_out_source786 = spike_out_source_array[786];
    end
    always @(spike_out_source_array[787]) begin 
        spike_out_source787 = spike_out_source_array[787];
    end
    always @(spike_out_source_array[788]) begin 
        spike_out_source788 = spike_out_source_array[788];
    end
    always @(spike_out_source_array[789]) begin 
        spike_out_source789 = spike_out_source_array[789];
    end
    always @(spike_out_source_array[790]) begin 
        spike_out_source790 = spike_out_source_array[790];
    end
    always @(spike_out_source_array[791]) begin 
        spike_out_source791 = spike_out_source_array[791];
    end
    always @(spike_out_source_array[792]) begin 
        spike_out_source792 = spike_out_source_array[792];
    end
    always @(spike_out_source_array[793]) begin 
        spike_out_source793 = spike_out_source_array[793];
    end
    always @(spike_out_source_array[794]) begin 
        spike_out_source794 = spike_out_source_array[794];
    end
    always @(spike_out_source_array[795]) begin 
        spike_out_source795 = spike_out_source_array[795];
    end
    always @(spike_out_source_array[796]) begin 
        spike_out_source796 = spike_out_source_array[796];
    end
    always @(spike_out_source_array[797]) begin 
        spike_out_source797 = spike_out_source_array[797];
    end
    always @(spike_out_source_array[798]) begin 
        spike_out_source798 = spike_out_source_array[798];
    end
    always @(spike_out_source_array[799]) begin 
        spike_out_source799 = spike_out_source_array[799];
    end
    always @(spike_out_source_array[800]) begin 
        spike_out_source800 = spike_out_source_array[800];
    end
    always @(spike_out_source_array[801]) begin 
        spike_out_source801 = spike_out_source_array[801];
    end
    always @(spike_out_source_array[802]) begin 
        spike_out_source802 = spike_out_source_array[802];
    end
    always @(spike_out_source_array[803]) begin 
        spike_out_source803 = spike_out_source_array[803];
    end
    always @(spike_out_source_array[804]) begin 
        spike_out_source804 = spike_out_source_array[804];
    end
    always @(spike_out_source_array[805]) begin 
        spike_out_source805 = spike_out_source_array[805];
    end
    always @(spike_out_source_array[806]) begin 
        spike_out_source806 = spike_out_source_array[806];
    end
    always @(spike_out_source_array[807]) begin 
        spike_out_source807 = spike_out_source_array[807];
    end
    always @(spike_out_source_array[808]) begin 
        spike_out_source808 = spike_out_source_array[808];
    end
    always @(spike_out_source_array[809]) begin 
        spike_out_source809 = spike_out_source_array[809];
    end
    always @(spike_out_source_array[810]) begin 
        spike_out_source810 = spike_out_source_array[810];
    end
    always @(spike_out_source_array[811]) begin 
        spike_out_source811 = spike_out_source_array[811];
    end
    always @(spike_out_source_array[812]) begin 
        spike_out_source812 = spike_out_source_array[812];
    end
    always @(spike_out_source_array[813]) begin 
        spike_out_source813 = spike_out_source_array[813];
    end
    always @(spike_out_source_array[814]) begin 
        spike_out_source814 = spike_out_source_array[814];
    end
    always @(spike_out_source_array[815]) begin 
        spike_out_source815 = spike_out_source_array[815];
    end
    always @(spike_out_source_array[816]) begin 
        spike_out_source816 = spike_out_source_array[816];
    end
    always @(spike_out_source_array[817]) begin 
        spike_out_source817 = spike_out_source_array[817];
    end
    always @(spike_out_source_array[818]) begin 
        spike_out_source818 = spike_out_source_array[818];
    end
    always @(spike_out_source_array[819]) begin 
        spike_out_source819 = spike_out_source_array[819];
    end
    always @(spike_out_source_array[820]) begin 
        spike_out_source820 = spike_out_source_array[820];
    end
    always @(spike_out_source_array[821]) begin 
        spike_out_source821 = spike_out_source_array[821];
    end
    always @(spike_out_source_array[822]) begin 
        spike_out_source822 = spike_out_source_array[822];
    end
    always @(spike_out_source_array[823]) begin 
        spike_out_source823 = spike_out_source_array[823];
    end
    always @(spike_out_source_array[824]) begin 
        spike_out_source824 = spike_out_source_array[824];
    end
    always @(spike_out_source_array[825]) begin 
        spike_out_source825 = spike_out_source_array[825];
    end
    always @(spike_out_source_array[826]) begin 
        spike_out_source826 = spike_out_source_array[826];
    end
    always @(spike_out_source_array[827]) begin 
        spike_out_source827 = spike_out_source_array[827];
    end
    always @(spike_out_source_array[828]) begin 
        spike_out_source828 = spike_out_source_array[828];
    end
    always @(spike_out_source_array[829]) begin 
        spike_out_source829 = spike_out_source_array[829];
    end
    always @(spike_out_source_array[830]) begin 
        spike_out_source830 = spike_out_source_array[830];
    end
    always @(spike_out_source_array[831]) begin 
        spike_out_source831 = spike_out_source_array[831];
    end
    always @(spike_out_source_array[832]) begin 
        spike_out_source832 = spike_out_source_array[832];
    end
    always @(spike_out_source_array[833]) begin 
        spike_out_source833 = spike_out_source_array[833];
    end
    always @(spike_out_source_array[834]) begin 
        spike_out_source834 = spike_out_source_array[834];
    end
    always @(spike_out_source_array[835]) begin 
        spike_out_source835 = spike_out_source_array[835];
    end
    always @(spike_out_source_array[836]) begin 
        spike_out_source836 = spike_out_source_array[836];
    end
    always @(spike_out_source_array[837]) begin 
        spike_out_source837 = spike_out_source_array[837];
    end
    always @(spike_out_source_array[838]) begin 
        spike_out_source838 = spike_out_source_array[838];
    end
    always @(spike_out_source_array[839]) begin 
        spike_out_source839 = spike_out_source_array[839];
    end
    always @(spike_out_source_array[840]) begin 
        spike_out_source840 = spike_out_source_array[840];
    end
    always @(spike_out_source_array[841]) begin 
        spike_out_source841 = spike_out_source_array[841];
    end
    always @(spike_out_source_array[842]) begin 
        spike_out_source842 = spike_out_source_array[842];
    end
    always @(spike_out_source_array[843]) begin 
        spike_out_source843 = spike_out_source_array[843];
    end
    always @(spike_out_source_array[844]) begin 
        spike_out_source844 = spike_out_source_array[844];
    end
    always @(spike_out_source_array[845]) begin 
        spike_out_source845 = spike_out_source_array[845];
    end
    always @(spike_out_source_array[846]) begin 
        spike_out_source846 = spike_out_source_array[846];
    end
    always @(spike_out_source_array[847]) begin 
        spike_out_source847 = spike_out_source_array[847];
    end
    always @(spike_out_source_array[848]) begin 
        spike_out_source848 = spike_out_source_array[848];
    end
    always @(spike_out_source_array[849]) begin 
        spike_out_source849 = spike_out_source_array[849];
    end
    always @(spike_out_source_array[850]) begin 
        spike_out_source850 = spike_out_source_array[850];
    end
    always @(spike_out_source_array[851]) begin 
        spike_out_source851 = spike_out_source_array[851];
    end
    always @(spike_out_source_array[852]) begin 
        spike_out_source852 = spike_out_source_array[852];
    end
    always @(spike_out_source_array[853]) begin 
        spike_out_source853 = spike_out_source_array[853];
    end
    always @(spike_out_source_array[854]) begin 
        spike_out_source854 = spike_out_source_array[854];
    end
    always @(spike_out_source_array[855]) begin 
        spike_out_source855 = spike_out_source_array[855];
    end
    always @(spike_out_source_array[856]) begin 
        spike_out_source856 = spike_out_source_array[856];
    end
    always @(spike_out_source_array[857]) begin 
        spike_out_source857 = spike_out_source_array[857];
    end
    always @(spike_out_source_array[858]) begin 
        spike_out_source858 = spike_out_source_array[858];
    end
    always @(spike_out_source_array[859]) begin 
        spike_out_source859 = spike_out_source_array[859];
    end
    always @(spike_out_source_array[860]) begin 
        spike_out_source860 = spike_out_source_array[860];
    end
    always @(spike_out_source_array[861]) begin 
        spike_out_source861 = spike_out_source_array[861];
    end
    always @(spike_out_source_array[862]) begin 
        spike_out_source862 = spike_out_source_array[862];
    end
    always @(spike_out_source_array[863]) begin 
        spike_out_source863 = spike_out_source_array[863];
    end
    always @(spike_out_source_array[864]) begin 
        spike_out_source864 = spike_out_source_array[864];
    end
    always @(spike_out_source_array[865]) begin 
        spike_out_source865 = spike_out_source_array[865];
    end
    always @(spike_out_source_array[866]) begin 
        spike_out_source866 = spike_out_source_array[866];
    end
    always @(spike_out_source_array[867]) begin 
        spike_out_source867 = spike_out_source_array[867];
    end
    always @(spike_out_source_array[868]) begin 
        spike_out_source868 = spike_out_source_array[868];
    end
    always @(spike_out_source_array[869]) begin 
        spike_out_source869 = spike_out_source_array[869];
    end
    always @(spike_out_source_array[870]) begin 
        spike_out_source870 = spike_out_source_array[870];
    end
    always @(spike_out_source_array[871]) begin 
        spike_out_source871 = spike_out_source_array[871];
    end
    always @(spike_out_source_array[872]) begin 
        spike_out_source872 = spike_out_source_array[872];
    end
    always @(spike_out_source_array[873]) begin 
        spike_out_source873 = spike_out_source_array[873];
    end
    always @(spike_out_source_array[874]) begin 
        spike_out_source874 = spike_out_source_array[874];
    end
    always @(spike_out_source_array[875]) begin 
        spike_out_source875 = spike_out_source_array[875];
    end
    always @(spike_out_source_array[876]) begin 
        spike_out_source876 = spike_out_source_array[876];
    end
    always @(spike_out_source_array[877]) begin 
        spike_out_source877 = spike_out_source_array[877];
    end
    always @(spike_out_source_array[878]) begin 
        spike_out_source878 = spike_out_source_array[878];
    end
    always @(spike_out_source_array[879]) begin 
        spike_out_source879 = spike_out_source_array[879];
    end
    always @(spike_out_source_array[880]) begin 
        spike_out_source880 = spike_out_source_array[880];
    end
    always @(spike_out_source_array[881]) begin 
        spike_out_source881 = spike_out_source_array[881];
    end
    always @(spike_out_source_array[882]) begin 
        spike_out_source882 = spike_out_source_array[882];
    end
    always @(spike_out_source_array[883]) begin 
        spike_out_source883 = spike_out_source_array[883];
    end
    always @(spike_out_source_array[884]) begin 
        spike_out_source884 = spike_out_source_array[884];
    end
    always @(spike_out_source_array[885]) begin 
        spike_out_source885 = spike_out_source_array[885];
    end
    always @(spike_out_source_array[886]) begin 
        spike_out_source886 = spike_out_source_array[886];
    end
    always @(spike_out_source_array[887]) begin 
        spike_out_source887 = spike_out_source_array[887];
    end
    always @(spike_out_source_array[888]) begin 
        spike_out_source888 = spike_out_source_array[888];
    end
    always @(spike_out_source_array[889]) begin 
        spike_out_source889 = spike_out_source_array[889];
    end
    always @(spike_out_source_array[890]) begin 
        spike_out_source890 = spike_out_source_array[890];
    end
    always @(spike_out_source_array[891]) begin 
        spike_out_source891 = spike_out_source_array[891];
    end
    always @(spike_out_source_array[892]) begin 
        spike_out_source892 = spike_out_source_array[892];
    end
    always @(spike_out_source_array[893]) begin 
        spike_out_source893 = spike_out_source_array[893];
    end
    always @(spike_out_source_array[894]) begin 
        spike_out_source894 = spike_out_source_array[894];
    end
    always @(spike_out_source_array[895]) begin 
        spike_out_source895 = spike_out_source_array[895];
    end
    always @(spike_out_source_array[896]) begin 
        spike_out_source896 = spike_out_source_array[896];
    end
    always @(spike_out_source_array[897]) begin 
        spike_out_source897 = spike_out_source_array[897];
    end
    always @(spike_out_source_array[898]) begin 
        spike_out_source898 = spike_out_source_array[898];
    end
    always @(spike_out_source_array[899]) begin 
        spike_out_source899 = spike_out_source_array[899];
    end
    always @(spike_out_source_array[900]) begin 
        spike_out_source900 = spike_out_source_array[900];
    end
    always @(spike_out_source_array[901]) begin 
        spike_out_source901 = spike_out_source_array[901];
    end
    always @(spike_out_source_array[902]) begin 
        spike_out_source902 = spike_out_source_array[902];
    end
    always @(spike_out_source_array[903]) begin 
        spike_out_source903 = spike_out_source_array[903];
    end
    always @(spike_out_source_array[904]) begin 
        spike_out_source904 = spike_out_source_array[904];
    end
    always @(spike_out_source_array[905]) begin 
        spike_out_source905 = spike_out_source_array[905];
    end
    always @(spike_out_source_array[906]) begin 
        spike_out_source906 = spike_out_source_array[906];
    end
    always @(spike_out_source_array[907]) begin 
        spike_out_source907 = spike_out_source_array[907];
    end
    always @(spike_out_source_array[908]) begin 
        spike_out_source908 = spike_out_source_array[908];
    end
    always @(spike_out_source_array[909]) begin 
        spike_out_source909 = spike_out_source_array[909];
    end
    always @(spike_out_source_array[910]) begin 
        spike_out_source910 = spike_out_source_array[910];
    end
    always @(spike_out_source_array[911]) begin 
        spike_out_source911 = spike_out_source_array[911];
    end
    always @(spike_out_source_array[912]) begin 
        spike_out_source912 = spike_out_source_array[912];
    end
    always @(spike_out_source_array[913]) begin 
        spike_out_source913 = spike_out_source_array[913];
    end
    always @(spike_out_source_array[914]) begin 
        spike_out_source914 = spike_out_source_array[914];
    end
    always @(spike_out_source_array[915]) begin 
        spike_out_source915 = spike_out_source_array[915];
    end
    always @(spike_out_source_array[916]) begin 
        spike_out_source916 = spike_out_source_array[916];
    end
    always @(spike_out_source_array[917]) begin 
        spike_out_source917 = spike_out_source_array[917];
    end
    always @(spike_out_source_array[918]) begin 
        spike_out_source918 = spike_out_source_array[918];
    end
    always @(spike_out_source_array[919]) begin 
        spike_out_source919 = spike_out_source_array[919];
    end
    always @(spike_out_source_array[920]) begin 
        spike_out_source920 = spike_out_source_array[920];
    end
    always @(spike_out_source_array[921]) begin 
        spike_out_source921 = spike_out_source_array[921];
    end
    always @(spike_out_source_array[922]) begin 
        spike_out_source922 = spike_out_source_array[922];
    end
    always @(spike_out_source_array[923]) begin 
        spike_out_source923 = spike_out_source_array[923];
    end
    always @(spike_out_source_array[924]) begin 
        spike_out_source924 = spike_out_source_array[924];
    end
    always @(spike_out_source_array[925]) begin 
        spike_out_source925 = spike_out_source_array[925];
    end
    always @(spike_out_source_array[926]) begin 
        spike_out_source926 = spike_out_source_array[926];
    end
    always @(spike_out_source_array[927]) begin 
        spike_out_source927 = spike_out_source_array[927];
    end
    always @(spike_out_source_array[928]) begin 
        spike_out_source928 = spike_out_source_array[928];
    end
    always @(spike_out_source_array[929]) begin 
        spike_out_source929 = spike_out_source_array[929];
    end
    always @(spike_out_source_array[930]) begin 
        spike_out_source930 = spike_out_source_array[930];
    end
    always @(spike_out_source_array[931]) begin 
        spike_out_source931 = spike_out_source_array[931];
    end
    always @(spike_out_source_array[932]) begin 
        spike_out_source932 = spike_out_source_array[932];
    end
    always @(spike_out_source_array[933]) begin 
        spike_out_source933 = spike_out_source_array[933];
    end
    always @(spike_out_source_array[934]) begin 
        spike_out_source934 = spike_out_source_array[934];
    end
    always @(spike_out_source_array[935]) begin 
        spike_out_source935 = spike_out_source_array[935];
    end
    always @(spike_out_source_array[936]) begin 
        spike_out_source936 = spike_out_source_array[936];
    end
    always @(spike_out_source_array[937]) begin 
        spike_out_source937 = spike_out_source_array[937];
    end
    always @(spike_out_source_array[938]) begin 
        spike_out_source938 = spike_out_source_array[938];
    end
    always @(spike_out_source_array[939]) begin 
        spike_out_source939 = spike_out_source_array[939];
    end
    always @(spike_out_source_array[940]) begin 
        spike_out_source940 = spike_out_source_array[940];
    end
    always @(spike_out_source_array[941]) begin 
        spike_out_source941 = spike_out_source_array[941];
    end
    always @(spike_out_source_array[942]) begin 
        spike_out_source942 = spike_out_source_array[942];
    end
    always @(spike_out_source_array[943]) begin 
        spike_out_source943 = spike_out_source_array[943];
    end
    always @(spike_out_source_array[944]) begin 
        spike_out_source944 = spike_out_source_array[944];
    end
    always @(spike_out_source_array[945]) begin 
        spike_out_source945 = spike_out_source_array[945];
    end
    always @(spike_out_source_array[946]) begin 
        spike_out_source946 = spike_out_source_array[946];
    end
    always @(spike_out_source_array[947]) begin 
        spike_out_source947 = spike_out_source_array[947];
    end
    always @(spike_out_source_array[948]) begin 
        spike_out_source948 = spike_out_source_array[948];
    end
    always @(spike_out_source_array[949]) begin 
        spike_out_source949 = spike_out_source_array[949];
    end
    always @(spike_out_source_array[950]) begin 
        spike_out_source950 = spike_out_source_array[950];
    end
    always @(spike_out_source_array[951]) begin 
        spike_out_source951 = spike_out_source_array[951];
    end
    always @(spike_out_source_array[952]) begin 
        spike_out_source952 = spike_out_source_array[952];
    end
    always @(spike_out_source_array[953]) begin 
        spike_out_source953 = spike_out_source_array[953];
    end
    always @(spike_out_source_array[954]) begin 
        spike_out_source954 = spike_out_source_array[954];
    end
    always @(spike_out_source_array[955]) begin 
        spike_out_source955 = spike_out_source_array[955];
    end
    always @(spike_out_source_array[956]) begin 
        spike_out_source956 = spike_out_source_array[956];
    end
    always @(spike_out_source_array[957]) begin 
        spike_out_source957 = spike_out_source_array[957];
    end
    always @(spike_out_source_array[958]) begin 
        spike_out_source958 = spike_out_source_array[958];
    end
    always @(spike_out_source_array[959]) begin 
        spike_out_source959 = spike_out_source_array[959];
    end
    always @(spike_out_source_array[960]) begin 
        spike_out_source960 = spike_out_source_array[960];
    end
    always @(spike_out_source_array[961]) begin 
        spike_out_source961 = spike_out_source_array[961];
    end
    always @(spike_out_source_array[962]) begin 
        spike_out_source962 = spike_out_source_array[962];
    end
    always @(spike_out_source_array[963]) begin 
        spike_out_source963 = spike_out_source_array[963];
    end
    always @(spike_out_source_array[964]) begin 
        spike_out_source964 = spike_out_source_array[964];
    end
    always @(spike_out_source_array[965]) begin 
        spike_out_source965 = spike_out_source_array[965];
    end
    always @(spike_out_source_array[966]) begin 
        spike_out_source966 = spike_out_source_array[966];
    end
    always @(spike_out_source_array[967]) begin 
        spike_out_source967 = spike_out_source_array[967];
    end
    always @(spike_out_source_array[968]) begin 
        spike_out_source968 = spike_out_source_array[968];
    end
    always @(spike_out_source_array[969]) begin 
        spike_out_source969 = spike_out_source_array[969];
    end
    always @(spike_out_source_array[970]) begin 
        spike_out_source970 = spike_out_source_array[970];
    end
    always @(spike_out_source_array[971]) begin 
        spike_out_source971 = spike_out_source_array[971];
    end
    always @(spike_out_source_array[972]) begin 
        spike_out_source972 = spike_out_source_array[972];
    end
    always @(spike_out_source_array[973]) begin 
        spike_out_source973 = spike_out_source_array[973];
    end
    always @(spike_out_source_array[974]) begin 
        spike_out_source974 = spike_out_source_array[974];
    end
    always @(spike_out_source_array[975]) begin 
        spike_out_source975 = spike_out_source_array[975];
    end
    always @(spike_out_source_array[976]) begin 
        spike_out_source976 = spike_out_source_array[976];
    end
    always @(spike_out_source_array[977]) begin 
        spike_out_source977 = spike_out_source_array[977];
    end
    always @(spike_out_source_array[978]) begin 
        spike_out_source978 = spike_out_source_array[978];
    end
    always @(spike_out_source_array[979]) begin 
        spike_out_source979 = spike_out_source_array[979];
    end
    always @(spike_out_source_array[980]) begin 
        spike_out_source980 = spike_out_source_array[980];
    end
    always @(spike_out_source_array[981]) begin 
        spike_out_source981 = spike_out_source_array[981];
    end
    always @(spike_out_source_array[982]) begin 
        spike_out_source982 = spike_out_source_array[982];
    end
    always @(spike_out_source_array[983]) begin 
        spike_out_source983 = spike_out_source_array[983];
    end
    always @(spike_out_source_array[984]) begin 
        spike_out_source984 = spike_out_source_array[984];
    end
    always @(spike_out_source_array[985]) begin 
        spike_out_source985 = spike_out_source_array[985];
    end
    always @(spike_out_source_array[986]) begin 
        spike_out_source986 = spike_out_source_array[986];
    end
    always @(spike_out_source_array[987]) begin 
        spike_out_source987 = spike_out_source_array[987];
    end
    always @(spike_out_source_array[988]) begin 
        spike_out_source988 = spike_out_source_array[988];
    end
    always @(spike_out_source_array[989]) begin 
        spike_out_source989 = spike_out_source_array[989];
    end
    always @(spike_out_source_array[990]) begin 
        spike_out_source990 = spike_out_source_array[990];
    end
    always @(spike_out_source_array[991]) begin 
        spike_out_source991 = spike_out_source_array[991];
    end
    always @(spike_out_source_array[992]) begin 
        spike_out_source992 = spike_out_source_array[992];
    end
    always @(spike_out_source_array[993]) begin 
        spike_out_source993 = spike_out_source_array[993];
    end
    always @(spike_out_source_array[994]) begin 
        spike_out_source994 = spike_out_source_array[994];
    end
    always @(spike_out_source_array[995]) begin 
        spike_out_source995 = spike_out_source_array[995];
    end
    always @(spike_out_source_array[996]) begin 
        spike_out_source996 = spike_out_source_array[996];
    end
    always @(spike_out_source_array[997]) begin 
        spike_out_source997 = spike_out_source_array[997];
    end
    always @(spike_out_source_array[998]) begin 
        spike_out_source998 = spike_out_source_array[998];
    end
    always @(spike_out_source_array[999]) begin 
        spike_out_source999 = spike_out_source_array[999];
    end
    always @(spike_out_source_array[1000]) begin 
        spike_out_source1000 = spike_out_source_array[1000];
    end
    always @(spike_out_source_array[1001]) begin 
        spike_out_source1001 = spike_out_source_array[1001];
    end
    always @(spike_out_source_array[1002]) begin 
        spike_out_source1002 = spike_out_source_array[1002];
    end
    always @(spike_out_source_array[1003]) begin 
        spike_out_source1003 = spike_out_source_array[1003];
    end
    always @(spike_out_source_array[1004]) begin 
        spike_out_source1004 = spike_out_source_array[1004];
    end
    always @(spike_out_source_array[1005]) begin 
        spike_out_source1005 = spike_out_source_array[1005];
    end
    always @(spike_out_source_array[1006]) begin 
        spike_out_source1006 = spike_out_source_array[1006];
    end
    always @(spike_out_source_array[1007]) begin 
        spike_out_source1007 = spike_out_source_array[1007];
    end
    always @(spike_out_source_array[1008]) begin 
        spike_out_source1008 = spike_out_source_array[1008];
    end
    always @(spike_out_source_array[1009]) begin 
        spike_out_source1009 = spike_out_source_array[1009];
    end
    always @(spike_out_source_array[1010]) begin 
        spike_out_source1010 = spike_out_source_array[1010];
    end
    always @(spike_out_source_array[1011]) begin 
        spike_out_source1011 = spike_out_source_array[1011];
    end
    always @(spike_out_source_array[1012]) begin 
        spike_out_source1012 = spike_out_source_array[1012];
    end
    always @(spike_out_source_array[1013]) begin 
        spike_out_source1013 = spike_out_source_array[1013];
    end
    always @(spike_out_source_array[1014]) begin 
        spike_out_source1014 = spike_out_source_array[1014];
    end
    always @(spike_out_source_array[1015]) begin 
        spike_out_source1015 = spike_out_source_array[1015];
    end
    always @(spike_out_source_array[1016]) begin 
        spike_out_source1016 = spike_out_source_array[1016];
    end
    always @(spike_out_source_array[1017]) begin 
        spike_out_source1017 = spike_out_source_array[1017];
    end
    always @(spike_out_source_array[1018]) begin 
        spike_out_source1018 = spike_out_source_array[1018];
    end
    always @(spike_out_source_array[1019]) begin 
        spike_out_source1019 = spike_out_source_array[1019];
    end
    always @(spike_out_source_array[1020]) begin 
        spike_out_source1020 = spike_out_source_array[1020];
    end
    always @(spike_out_source_array[1021]) begin 
        spike_out_source1021 = spike_out_source_array[1021];
    end
    always @(spike_out_source_array[1022]) begin 
        spike_out_source1022 = spike_out_source_array[1022];
    end
    always @(spike_out_source_array[1023]) begin 
        spike_out_source1023 = spike_out_source_array[1023];
    end
    reg[18:0] i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21;
    reg[18:0] j1, j2, j3, j4, j5, j6, j7, j8, j9, j10, j11, j12, j13, j14, j15, j16, j17, j18, j19, j20, j21;
    network_interface_scaled ni1(
        .spike_out_source0(spike_out_source[0]),
        .spike_out_source1(spike_out_source[1]),        .spike_out_source2(spike_out_source[2]),        .spike_out_source3(spike_out_source[3]),        .spike_out_source4(spike_out_source[4]),        .spike_out_source5(spike_out_source[5]),        .spike_out_source6(spike_out_source[6]),        .spike_out_source7(spike_out_source[7]),        .spike_out_source8(spike_out_source[8]),        .spike_out_source9(spike_out_source[9]),        .spike_out_source10(spike_out_source[10]),        .spike_out_source11(spike_out_source[11]),        .spike_out_source12(spike_out_source[12]),        .spike_out_source13(spike_out_source[13]),        .spike_out_source14(spike_out_source[14]),        .spike_out_source15(spike_out_source[15]),        .spike_out_source16(spike_out_source[16]),        .spike_out_source17(spike_out_source[17]),        .spike_out_source18(spike_out_source[18]),        .spike_out_source19(spike_out_source[19]),        .spike_out_source20(spike_out_source[20]),        .spike_out_source21(spike_out_source[21]),        .spike_out_source22(spike_out_source[22]),        .spike_out_source23(spike_out_source[23]),        .spike_out_source24(spike_out_source[24]),        .spike_out_source25(spike_out_source[25]),        .spike_out_source26(spike_out_source[26]),        .spike_out_source27(spike_out_source[27]),        .spike_out_source28(spike_out_source[28]),        .spike_out_source29(spike_out_source[29]),        .spike_out_source30(spike_out_source[30]),        .spike_out_source31(spike_out_source[31]),        .spike_out_source32(spike_out_source[32]),        .spike_out_source33(spike_out_source[33]),        .spike_out_source34(spike_out_source[34]),        .spike_out_source35(spike_out_source[35]),        .spike_out_source36(spike_out_source[36]),        .spike_out_source37(spike_out_source[37]),        .spike_out_source38(spike_out_source[38]),        .spike_out_source39(spike_out_source[39]),        .spike_out_source40(spike_out_source[40]),        .spike_out_source41(spike_out_source[41]),        .spike_out_source42(spike_out_source[42]),        .spike_out_source43(spike_out_source[43]),        .spike_out_source44(spike_out_source[44]),        .spike_out_source45(spike_out_source[45]),        .spike_out_source46(spike_out_source[46]),        .spike_out_source47(spike_out_source[47]),        .spike_out_source48(spike_out_source[48]),        .spike_out_source49(spike_out_source[49]),        .spike_out_source50(spike_out_source[50]),        .spike_out_source51(spike_out_source[51]),        .spike_out_source52(spike_out_source[52]),        .spike_out_source53(spike_out_source[53]),        .spike_out_source54(spike_out_source[54]),        .spike_out_source55(spike_out_source[55]),        .spike_out_source56(spike_out_source[56]),        .spike_out_source57(spike_out_source[57]),        .spike_out_source58(spike_out_source[58]),        .spike_out_source59(spike_out_source[59]),        .spike_out_source60(spike_out_source[60]),        .spike_out_source61(spike_out_source[61]),        .spike_out_source62(spike_out_source[62]),        .spike_out_source63(spike_out_source[63]),        .spike_out_source64(spike_out_source[64]),        .spike_out_source65(spike_out_source[65]),        .spike_out_source66(spike_out_source[66]),        .spike_out_source67(spike_out_source[67]),        .spike_out_source68(spike_out_source[68]),        .spike_out_source69(spike_out_source[69]),        .spike_out_source70(spike_out_source[70]),        .spike_out_source71(spike_out_source[71]),        .spike_out_source72(spike_out_source[72]),        .spike_out_source73(spike_out_source[73]),        .spike_out_source74(spike_out_source[74]),        .spike_out_source75(spike_out_source[75]),        .spike_out_source76(spike_out_source[76]),        .spike_out_source77(spike_out_source[77]),        .spike_out_source78(spike_out_source[78]),        .spike_out_source79(spike_out_source[79]),        .spike_out_source80(spike_out_source[80]),        .spike_out_source81(spike_out_source[81]),        .spike_out_source82(spike_out_source[82]),        .spike_out_source83(spike_out_source[83]),        .spike_out_source84(spike_out_source[84]),        .spike_out_source85(spike_out_source[85]),        .spike_out_source86(spike_out_source[86]),        .spike_out_source87(spike_out_source[87]),        .spike_out_source88(spike_out_source[88]),        .spike_out_source89(spike_out_source[89]),        .spike_out_source90(spike_out_source[90]),        .spike_out_source91(spike_out_source[91]),        .spike_out_source92(spike_out_source[92]),        .spike_out_source93(spike_out_source[93]),        .spike_out_source94(spike_out_source[94]),        .spike_out_source95(spike_out_source[95]),        .spike_out_source96(spike_out_source[96]),        .spike_out_source97(spike_out_source[97]),        .spike_out_source98(spike_out_source[98]),        .spike_out_source99(spike_out_source[99]),        .spike_out_source100(spike_out_source[100]),
        .spike_out_source101(spike_out_source[101]),        .spike_out_source102(spike_out_source[102]),        .spike_out_source103(spike_out_source[103]),        .spike_out_source104(spike_out_source[104]),        .spike_out_source105(spike_out_source[105]),        .spike_out_source106(spike_out_source[106]),        .spike_out_source107(spike_out_source[107]),        .spike_out_source108(spike_out_source[108]),        .spike_out_source109(spike_out_source[109]),        .spike_out_source110(spike_out_source[110]),        .spike_out_source111(spike_out_source[111]),        .spike_out_source112(spike_out_source[112]),        .spike_out_source113(spike_out_source[113]),        .spike_out_source114(spike_out_source[114]),        .spike_out_source115(spike_out_source[115]),        .spike_out_source116(spike_out_source[116]),        .spike_out_source117(spike_out_source[117]),        .spike_out_source118(spike_out_source[118]),        .spike_out_source119(spike_out_source[119]),        .spike_out_source120(spike_out_source[120]),        .spike_out_source121(spike_out_source[121]),        .spike_out_source122(spike_out_source[122]),        .spike_out_source123(spike_out_source[123]),        .spike_out_source124(spike_out_source[124]),        .spike_out_source125(spike_out_source[125]),        .spike_out_source126(spike_out_source[126]),        .spike_out_source127(spike_out_source[127]),        .spike_out_source128(spike_out_source[128]),        .spike_out_source129(spike_out_source[129]),        .spike_out_source130(spike_out_source[130]),        .spike_out_source131(spike_out_source[131]),        .spike_out_source132(spike_out_source[132]),        .spike_out_source133(spike_out_source[133]),        .spike_out_source134(spike_out_source[134]),        .spike_out_source135(spike_out_source[135]),        .spike_out_source136(spike_out_source[136]),        .spike_out_source137(spike_out_source[137]),        .spike_out_source138(spike_out_source[138]),        .spike_out_source139(spike_out_source[139]),        .spike_out_source140(spike_out_source[140]),        .spike_out_source141(spike_out_source[141]),        .spike_out_source142(spike_out_source[142]),        .spike_out_source143(spike_out_source[143]),        .spike_out_source144(spike_out_source[144]),        .spike_out_source145(spike_out_source[145]),        .spike_out_source146(spike_out_source[146]),        .spike_out_source147(spike_out_source[147]),        .spike_out_source148(spike_out_source[148]),        .spike_out_source149(spike_out_source[149]),        .spike_out_source150(spike_out_source[150]),        .spike_out_source151(spike_out_source[151]),        .spike_out_source152(spike_out_source[152]),        .spike_out_source153(spike_out_source[153]),        .spike_out_source154(spike_out_source[154]),        .spike_out_source155(spike_out_source[155]),        .spike_out_source156(spike_out_source[156]),        .spike_out_source157(spike_out_source[157]),        .spike_out_source158(spike_out_source[158]),        .spike_out_source159(spike_out_source[159]),        .spike_out_source160(spike_out_source[160]),        .spike_out_source161(spike_out_source[161]),        .spike_out_source162(spike_out_source[162]),        .spike_out_source163(spike_out_source[163]),        .spike_out_source164(spike_out_source[164]),        .spike_out_source165(spike_out_source[165]),        .spike_out_source166(spike_out_source[166]),        .spike_out_source167(spike_out_source[167]),        .spike_out_source168(spike_out_source[168]),        .spike_out_source169(spike_out_source[169]),        .spike_out_source170(spike_out_source[170]),        .spike_out_source171(spike_out_source[171]),        .spike_out_source172(spike_out_source[172]),        .spike_out_source173(spike_out_source[173]),        .spike_out_source174(spike_out_source[174]),        .spike_out_source175(spike_out_source[175]),        .spike_out_source176(spike_out_source[176]),        .spike_out_source177(spike_out_source[177]),        .spike_out_source178(spike_out_source[178]),        .spike_out_source179(spike_out_source[179]),        .spike_out_source180(spike_out_source[180]),        .spike_out_source181(spike_out_source[181]),        .spike_out_source182(spike_out_source[182]),        .spike_out_source183(spike_out_source[183]),        .spike_out_source184(spike_out_source[184]),        .spike_out_source185(spike_out_source[185]),        .spike_out_source186(spike_out_source[186]),        .spike_out_source187(spike_out_source[187]),        .spike_out_source188(spike_out_source[188]),        .spike_out_source189(spike_out_source[189]),        .spike_out_source190(spike_out_source[190]),        .spike_out_source191(spike_out_source[191]),        .spike_out_source192(spike_out_source[192]),        .spike_out_source193(spike_out_source[193]),        .spike_out_source194(spike_out_source[194]),        .spike_out_source195(spike_out_source[195]),        .spike_out_source196(spike_out_source[196]),        .spike_out_source197(spike_out_source[197]),        .spike_out_source198(spike_out_source[198]),        .spike_out_source199(spike_out_source[199]),        .spike_out_source200(spike_out_source[200]),
        .spike_out_source201(spike_out_source[201]),        .spike_out_source202(spike_out_source[202]),        .spike_out_source203(spike_out_source[203]),        .spike_out_source204(spike_out_source[204]),        .spike_out_source205(spike_out_source[205]),        .spike_out_source206(spike_out_source[206]),        .spike_out_source207(spike_out_source[207]),        .spike_out_source208(spike_out_source[208]),        .spike_out_source209(spike_out_source[209]),        .spike_out_source210(spike_out_source[210]),        .spike_out_source211(spike_out_source[211]),        .spike_out_source212(spike_out_source[212]),        .spike_out_source213(spike_out_source[213]),        .spike_out_source214(spike_out_source[214]),        .spike_out_source215(spike_out_source[215]),        .spike_out_source216(spike_out_source[216]),        .spike_out_source217(spike_out_source[217]),        .spike_out_source218(spike_out_source[218]),        .spike_out_source219(spike_out_source[219]),        .spike_out_source220(spike_out_source[220]),        .spike_out_source221(spike_out_source[221]),        .spike_out_source222(spike_out_source[222]),        .spike_out_source223(spike_out_source[223]),        .spike_out_source224(spike_out_source[224]),        .spike_out_source225(spike_out_source[225]),        .spike_out_source226(spike_out_source[226]),        .spike_out_source227(spike_out_source[227]),        .spike_out_source228(spike_out_source[228]),        .spike_out_source229(spike_out_source[229]),        .spike_out_source230(spike_out_source[230]),        .spike_out_source231(spike_out_source[231]),        .spike_out_source232(spike_out_source[232]),        .spike_out_source233(spike_out_source[233]),        .spike_out_source234(spike_out_source[234]),        .spike_out_source235(spike_out_source[235]),        .spike_out_source236(spike_out_source[236]),        .spike_out_source237(spike_out_source[237]),        .spike_out_source238(spike_out_source[238]),        .spike_out_source239(spike_out_source[239]),        .spike_out_source240(spike_out_source[240]),        .spike_out_source241(spike_out_source[241]),        .spike_out_source242(spike_out_source[242]),        .spike_out_source243(spike_out_source[243]),        .spike_out_source244(spike_out_source[244]),        .spike_out_source245(spike_out_source[245]),        .spike_out_source246(spike_out_source[246]),        .spike_out_source247(spike_out_source[247]),        .spike_out_source248(spike_out_source[248]),        .spike_out_source249(spike_out_source[249]),        .spike_out_source250(spike_out_source[250]),        .spike_out_source251(spike_out_source[251]),        .spike_out_source252(spike_out_source[252]),        .spike_out_source253(spike_out_source[253]),        .spike_out_source254(spike_out_source[254]),        .spike_out_source255(spike_out_source[255]),        .spike_out_source256(spike_out_source[256]),        .spike_out_source257(spike_out_source[257]),        .spike_out_source258(spike_out_source[258]),        .spike_out_source259(spike_out_source[259]),        .spike_out_source260(spike_out_source[260]),        .spike_out_source261(spike_out_source[261]),        .spike_out_source262(spike_out_source[262]),        .spike_out_source263(spike_out_source[263]),        .spike_out_source264(spike_out_source[264]),        .spike_out_source265(spike_out_source[265]),        .spike_out_source266(spike_out_source[266]),        .spike_out_source267(spike_out_source[267]),        .spike_out_source268(spike_out_source[268]),        .spike_out_source269(spike_out_source[269]),        .spike_out_source270(spike_out_source[270]),        .spike_out_source271(spike_out_source[271]),        .spike_out_source272(spike_out_source[272]),        .spike_out_source273(spike_out_source[273]),        .spike_out_source274(spike_out_source[274]),        .spike_out_source275(spike_out_source[275]),        .spike_out_source276(spike_out_source[276]),        .spike_out_source277(spike_out_source[277]),        .spike_out_source278(spike_out_source[278]),        .spike_out_source279(spike_out_source[279]),        .spike_out_source280(spike_out_source[280]),        .spike_out_source281(spike_out_source[281]),        .spike_out_source282(spike_out_source[282]),        .spike_out_source283(spike_out_source[283]),        .spike_out_source284(spike_out_source[284]),        .spike_out_source285(spike_out_source[285]),        .spike_out_source286(spike_out_source[286]),        .spike_out_source287(spike_out_source[287]),        .spike_out_source288(spike_out_source[288]),        .spike_out_source289(spike_out_source[289]),        .spike_out_source290(spike_out_source[290]),        .spike_out_source291(spike_out_source[291]),        .spike_out_source292(spike_out_source[292]),        .spike_out_source293(spike_out_source[293]),        .spike_out_source294(spike_out_source[294]),        .spike_out_source295(spike_out_source[295]),        .spike_out_source296(spike_out_source[296]),        .spike_out_source297(spike_out_source[297]),        .spike_out_source298(spike_out_source[298]),        .spike_out_source299(spike_out_source[299]),        .spike_out_source300(spike_out_source[300]),
        .spike_out_source301(spike_out_source[301]),        .spike_out_source302(spike_out_source[302]),        .spike_out_source303(spike_out_source[303]),        .spike_out_source304(spike_out_source[304]),        .spike_out_source305(spike_out_source[305]),        .spike_out_source306(spike_out_source[306]),        .spike_out_source307(spike_out_source[307]),        .spike_out_source308(spike_out_source[308]),        .spike_out_source309(spike_out_source[309]),        .spike_out_source310(spike_out_source[310]),        .spike_out_source311(spike_out_source[311]),        .spike_out_source312(spike_out_source[312]),        .spike_out_source313(spike_out_source[313]),        .spike_out_source314(spike_out_source[314]),        .spike_out_source315(spike_out_source[315]),        .spike_out_source316(spike_out_source[316]),        .spike_out_source317(spike_out_source[317]),        .spike_out_source318(spike_out_source[318]),        .spike_out_source319(spike_out_source[319]),        .spike_out_source320(spike_out_source[320]),        .spike_out_source321(spike_out_source[321]),        .spike_out_source322(spike_out_source[322]),        .spike_out_source323(spike_out_source[323]),        .spike_out_source324(spike_out_source[324]),        .spike_out_source325(spike_out_source[325]),        .spike_out_source326(spike_out_source[326]),        .spike_out_source327(spike_out_source[327]),        .spike_out_source328(spike_out_source[328]),        .spike_out_source329(spike_out_source[329]),        .spike_out_source330(spike_out_source[330]),        .spike_out_source331(spike_out_source[331]),        .spike_out_source332(spike_out_source[332]),        .spike_out_source333(spike_out_source[333]),        .spike_out_source334(spike_out_source[334]),        .spike_out_source335(spike_out_source[335]),        .spike_out_source336(spike_out_source[336]),        .spike_out_source337(spike_out_source[337]),        .spike_out_source338(spike_out_source[338]),        .spike_out_source339(spike_out_source[339]),        .spike_out_source340(spike_out_source[340]),        .spike_out_source341(spike_out_source[341]),        .spike_out_source342(spike_out_source[342]),        .spike_out_source343(spike_out_source[343]),        .spike_out_source344(spike_out_source[344]),        .spike_out_source345(spike_out_source[345]),        .spike_out_source346(spike_out_source[346]),        .spike_out_source347(spike_out_source[347]),        .spike_out_source348(spike_out_source[348]),        .spike_out_source349(spike_out_source[349]),        .spike_out_source350(spike_out_source[350]),        .spike_out_source351(spike_out_source[351]),        .spike_out_source352(spike_out_source[352]),        .spike_out_source353(spike_out_source[353]),        .spike_out_source354(spike_out_source[354]),        .spike_out_source355(spike_out_source[355]),        .spike_out_source356(spike_out_source[356]),        .spike_out_source357(spike_out_source[357]),        .spike_out_source358(spike_out_source[358]),        .spike_out_source359(spike_out_source[359]),        .spike_out_source360(spike_out_source[360]),        .spike_out_source361(spike_out_source[361]),        .spike_out_source362(spike_out_source[362]),        .spike_out_source363(spike_out_source[363]),        .spike_out_source364(spike_out_source[364]),        .spike_out_source365(spike_out_source[365]),        .spike_out_source366(spike_out_source[366]),        .spike_out_source367(spike_out_source[367]),        .spike_out_source368(spike_out_source[368]),        .spike_out_source369(spike_out_source[369]),        .spike_out_source370(spike_out_source[370]),        .spike_out_source371(spike_out_source[371]),        .spike_out_source372(spike_out_source[372]),        .spike_out_source373(spike_out_source[373]),        .spike_out_source374(spike_out_source[374]),        .spike_out_source375(spike_out_source[375]),        .spike_out_source376(spike_out_source[376]),        .spike_out_source377(spike_out_source[377]),        .spike_out_source378(spike_out_source[378]),        .spike_out_source379(spike_out_source[379]),        .spike_out_source380(spike_out_source[380]),        .spike_out_source381(spike_out_source[381]),        .spike_out_source382(spike_out_source[382]),        .spike_out_source383(spike_out_source[383]),        .spike_out_source384(spike_out_source[384]),        .spike_out_source385(spike_out_source[385]),        .spike_out_source386(spike_out_source[386]),        .spike_out_source387(spike_out_source[387]),        .spike_out_source388(spike_out_source[388]),        .spike_out_source389(spike_out_source[389]),        .spike_out_source390(spike_out_source[390]),        .spike_out_source391(spike_out_source[391]),        .spike_out_source392(spike_out_source[392]),        .spike_out_source393(spike_out_source[393]),        .spike_out_source394(spike_out_source[394]),        .spike_out_source395(spike_out_source[395]),        .spike_out_source396(spike_out_source[396]),        .spike_out_source397(spike_out_source[397]),        .spike_out_source398(spike_out_source[398]),        .spike_out_source399(spike_out_source[399]),        .spike_out_source400(spike_out_source[400]),
        .spike_out_source401(spike_out_source[401]),        .spike_out_source402(spike_out_source[402]),        .spike_out_source403(spike_out_source[403]),        .spike_out_source404(spike_out_source[404]),        .spike_out_source405(spike_out_source[405]),        .spike_out_source406(spike_out_source[406]),        .spike_out_source407(spike_out_source[407]),        .spike_out_source408(spike_out_source[408]),        .spike_out_source409(spike_out_source[409]),        .spike_out_source410(spike_out_source[410]),        .spike_out_source411(spike_out_source[411]),        .spike_out_source412(spike_out_source[412]),        .spike_out_source413(spike_out_source[413]),        .spike_out_source414(spike_out_source[414]),        .spike_out_source415(spike_out_source[415]),        .spike_out_source416(spike_out_source[416]),        .spike_out_source417(spike_out_source[417]),        .spike_out_source418(spike_out_source[418]),        .spike_out_source419(spike_out_source[419]),        .spike_out_source420(spike_out_source[420]),        .spike_out_source421(spike_out_source[421]),        .spike_out_source422(spike_out_source[422]),        .spike_out_source423(spike_out_source[423]),        .spike_out_source424(spike_out_source[424]),        .spike_out_source425(spike_out_source[425]),        .spike_out_source426(spike_out_source[426]),        .spike_out_source427(spike_out_source[427]),        .spike_out_source428(spike_out_source[428]),        .spike_out_source429(spike_out_source[429]),        .spike_out_source430(spike_out_source[430]),        .spike_out_source431(spike_out_source[431]),        .spike_out_source432(spike_out_source[432]),        .spike_out_source433(spike_out_source[433]),        .spike_out_source434(spike_out_source[434]),        .spike_out_source435(spike_out_source[435]),        .spike_out_source436(spike_out_source[436]),        .spike_out_source437(spike_out_source[437]),        .spike_out_source438(spike_out_source[438]),        .spike_out_source439(spike_out_source[439]),        .spike_out_source440(spike_out_source[440]),        .spike_out_source441(spike_out_source[441]),        .spike_out_source442(spike_out_source[442]),        .spike_out_source443(spike_out_source[443]),        .spike_out_source444(spike_out_source[444]),        .spike_out_source445(spike_out_source[445]),        .spike_out_source446(spike_out_source[446]),        .spike_out_source447(spike_out_source[447]),        .spike_out_source448(spike_out_source[448]),        .spike_out_source449(spike_out_source[449]),        .spike_out_source450(spike_out_source[450]),        .spike_out_source451(spike_out_source[451]),        .spike_out_source452(spike_out_source[452]),        .spike_out_source453(spike_out_source[453]),        .spike_out_source454(spike_out_source[454]),        .spike_out_source455(spike_out_source[455]),        .spike_out_source456(spike_out_source[456]),        .spike_out_source457(spike_out_source[457]),        .spike_out_source458(spike_out_source[458]),        .spike_out_source459(spike_out_source[459]),        .spike_out_source460(spike_out_source[460]),        .spike_out_source461(spike_out_source[461]),        .spike_out_source462(spike_out_source[462]),        .spike_out_source463(spike_out_source[463]),        .spike_out_source464(spike_out_source[464]),        .spike_out_source465(spike_out_source[465]),        .spike_out_source466(spike_out_source[466]),        .spike_out_source467(spike_out_source[467]),        .spike_out_source468(spike_out_source[468]),        .spike_out_source469(spike_out_source[469]),        .spike_out_source470(spike_out_source[470]),        .spike_out_source471(spike_out_source[471]),        .spike_out_source472(spike_out_source[472]),        .spike_out_source473(spike_out_source[473]),        .spike_out_source474(spike_out_source[474]),        .spike_out_source475(spike_out_source[475]),        .spike_out_source476(spike_out_source[476]),        .spike_out_source477(spike_out_source[477]),        .spike_out_source478(spike_out_source[478]),        .spike_out_source479(spike_out_source[479]),        .spike_out_source480(spike_out_source[480]),        .spike_out_source481(spike_out_source[481]),        .spike_out_source482(spike_out_source[482]),        .spike_out_source483(spike_out_source[483]),        .spike_out_source484(spike_out_source[484]),        .spike_out_source485(spike_out_source[485]),        .spike_out_source486(spike_out_source[486]),        .spike_out_source487(spike_out_source[487]),        .spike_out_source488(spike_out_source[488]),        .spike_out_source489(spike_out_source[489]),        .spike_out_source490(spike_out_source[490]),        .spike_out_source491(spike_out_source[491]),        .spike_out_source492(spike_out_source[492]),        .spike_out_source493(spike_out_source[493]),        .spike_out_source494(spike_out_source[494]),        .spike_out_source495(spike_out_source[495]),        .spike_out_source496(spike_out_source[496]),        .spike_out_source497(spike_out_source[497]),        .spike_out_source498(spike_out_source[498]),        .spike_out_source499(spike_out_source[499]),        .spike_out_source500(spike_out_source[500]),
        .spike_out_source501(spike_out_source[501]),        .spike_out_source502(spike_out_source[502]),        .spike_out_source503(spike_out_source[503]),        .spike_out_source504(spike_out_source[504]),        .spike_out_source505(spike_out_source[505]),        .spike_out_source506(spike_out_source[506]),        .spike_out_source507(spike_out_source[507]),        .spike_out_source508(spike_out_source[508]),        .spike_out_source509(spike_out_source[509]),        .spike_out_source510(spike_out_source[510]),        .spike_out_source511(spike_out_source[511]),        .spike_out_source512(spike_out_source[512]),        .spike_out_source513(spike_out_source[513]),        .spike_out_source514(spike_out_source[514]),        .spike_out_source515(spike_out_source[515]),        .spike_out_source516(spike_out_source[516]),        .spike_out_source517(spike_out_source[517]),        .spike_out_source518(spike_out_source[518]),        .spike_out_source519(spike_out_source[519]),        .spike_out_source520(spike_out_source[520]),        .spike_out_source521(spike_out_source[521]),        .spike_out_source522(spike_out_source[522]),        .spike_out_source523(spike_out_source[523]),        .spike_out_source524(spike_out_source[524]),        .spike_out_source525(spike_out_source[525]),        .spike_out_source526(spike_out_source[526]),        .spike_out_source527(spike_out_source[527]),        .spike_out_source528(spike_out_source[528]),        .spike_out_source529(spike_out_source[529]),        .spike_out_source530(spike_out_source[530]),        .spike_out_source531(spike_out_source[531]),        .spike_out_source532(spike_out_source[532]),        .spike_out_source533(spike_out_source[533]),        .spike_out_source534(spike_out_source[534]),        .spike_out_source535(spike_out_source[535]),        .spike_out_source536(spike_out_source[536]),        .spike_out_source537(spike_out_source[537]),        .spike_out_source538(spike_out_source[538]),        .spike_out_source539(spike_out_source[539]),        .spike_out_source540(spike_out_source[540]),        .spike_out_source541(spike_out_source[541]),        .spike_out_source542(spike_out_source[542]),        .spike_out_source543(spike_out_source[543]),        .spike_out_source544(spike_out_source[544]),        .spike_out_source545(spike_out_source[545]),        .spike_out_source546(spike_out_source[546]),        .spike_out_source547(spike_out_source[547]),        .spike_out_source548(spike_out_source[548]),        .spike_out_source549(spike_out_source[549]),        .spike_out_source550(spike_out_source[550]),        .spike_out_source551(spike_out_source[551]),        .spike_out_source552(spike_out_source[552]),        .spike_out_source553(spike_out_source[553]),        .spike_out_source554(spike_out_source[554]),        .spike_out_source555(spike_out_source[555]),        .spike_out_source556(spike_out_source[556]),        .spike_out_source557(spike_out_source[557]),        .spike_out_source558(spike_out_source[558]),        .spike_out_source559(spike_out_source[559]),        .spike_out_source560(spike_out_source[560]),        .spike_out_source561(spike_out_source[561]),        .spike_out_source562(spike_out_source[562]),        .spike_out_source563(spike_out_source[563]),        .spike_out_source564(spike_out_source[564]),        .spike_out_source565(spike_out_source[565]),        .spike_out_source566(spike_out_source[566]),        .spike_out_source567(spike_out_source[567]),        .spike_out_source568(spike_out_source[568]),        .spike_out_source569(spike_out_source[569]),        .spike_out_source570(spike_out_source[570]),        .spike_out_source571(spike_out_source[571]),        .spike_out_source572(spike_out_source[572]),        .spike_out_source573(spike_out_source[573]),        .spike_out_source574(spike_out_source[574]),        .spike_out_source575(spike_out_source[575]),        .spike_out_source576(spike_out_source[576]),        .spike_out_source577(spike_out_source[577]),        .spike_out_source578(spike_out_source[578]),        .spike_out_source579(spike_out_source[579]),        .spike_out_source580(spike_out_source[580]),        .spike_out_source581(spike_out_source[581]),        .spike_out_source582(spike_out_source[582]),        .spike_out_source583(spike_out_source[583]),        .spike_out_source584(spike_out_source[584]),        .spike_out_source585(spike_out_source[585]),        .spike_out_source586(spike_out_source[586]),        .spike_out_source587(spike_out_source[587]),        .spike_out_source588(spike_out_source[588]),        .spike_out_source589(spike_out_source[589]),        .spike_out_source590(spike_out_source[590]),        .spike_out_source591(spike_out_source[591]),        .spike_out_source592(spike_out_source[592]),        .spike_out_source593(spike_out_source[593]),        .spike_out_source594(spike_out_source[594]),        .spike_out_source595(spike_out_source[595]),        .spike_out_source596(spike_out_source[596]),        .spike_out_source597(spike_out_source[597]),        .spike_out_source598(spike_out_source[598]),        .spike_out_source599(spike_out_source[599]),        .spike_out_source600(spike_out_source[600]),
        .spike_out_source601(spike_out_source[601]),        .spike_out_source602(spike_out_source[602]),        .spike_out_source603(spike_out_source[603]),        .spike_out_source604(spike_out_source[604]),        .spike_out_source605(spike_out_source[605]),        .spike_out_source606(spike_out_source[606]),        .spike_out_source607(spike_out_source[607]),        .spike_out_source608(spike_out_source[608]),        .spike_out_source609(spike_out_source[609]),        .spike_out_source610(spike_out_source[610]),        .spike_out_source611(spike_out_source[611]),        .spike_out_source612(spike_out_source[612]),        .spike_out_source613(spike_out_source[613]),        .spike_out_source614(spike_out_source[614]),        .spike_out_source615(spike_out_source[615]),        .spike_out_source616(spike_out_source[616]),        .spike_out_source617(spike_out_source[617]),        .spike_out_source618(spike_out_source[618]),        .spike_out_source619(spike_out_source[619]),        .spike_out_source620(spike_out_source[620]),        .spike_out_source621(spike_out_source[621]),        .spike_out_source622(spike_out_source[622]),        .spike_out_source623(spike_out_source[623]),        .spike_out_source624(spike_out_source[624]),        .spike_out_source625(spike_out_source[625]),        .spike_out_source626(spike_out_source[626]),        .spike_out_source627(spike_out_source[627]),        .spike_out_source628(spike_out_source[628]),        .spike_out_source629(spike_out_source[629]),        .spike_out_source630(spike_out_source[630]),        .spike_out_source631(spike_out_source[631]),        .spike_out_source632(spike_out_source[632]),        .spike_out_source633(spike_out_source[633]),        .spike_out_source634(spike_out_source[634]),        .spike_out_source635(spike_out_source[635]),        .spike_out_source636(spike_out_source[636]),        .spike_out_source637(spike_out_source[637]),        .spike_out_source638(spike_out_source[638]),        .spike_out_source639(spike_out_source[639]),        .spike_out_source640(spike_out_source[640]),        .spike_out_source641(spike_out_source[641]),        .spike_out_source642(spike_out_source[642]),        .spike_out_source643(spike_out_source[643]),        .spike_out_source644(spike_out_source[644]),        .spike_out_source645(spike_out_source[645]),        .spike_out_source646(spike_out_source[646]),        .spike_out_source647(spike_out_source[647]),        .spike_out_source648(spike_out_source[648]),        .spike_out_source649(spike_out_source[649]),        .spike_out_source650(spike_out_source[650]),        .spike_out_source651(spike_out_source[651]),        .spike_out_source652(spike_out_source[652]),        .spike_out_source653(spike_out_source[653]),        .spike_out_source654(spike_out_source[654]),        .spike_out_source655(spike_out_source[655]),        .spike_out_source656(spike_out_source[656]),        .spike_out_source657(spike_out_source[657]),        .spike_out_source658(spike_out_source[658]),        .spike_out_source659(spike_out_source[659]),        .spike_out_source660(spike_out_source[660]),        .spike_out_source661(spike_out_source[661]),        .spike_out_source662(spike_out_source[662]),        .spike_out_source663(spike_out_source[663]),        .spike_out_source664(spike_out_source[664]),        .spike_out_source665(spike_out_source[665]),        .spike_out_source666(spike_out_source[666]),        .spike_out_source667(spike_out_source[667]),        .spike_out_source668(spike_out_source[668]),        .spike_out_source669(spike_out_source[669]),        .spike_out_source670(spike_out_source[670]),        .spike_out_source671(spike_out_source[671]),        .spike_out_source672(spike_out_source[672]),        .spike_out_source673(spike_out_source[673]),        .spike_out_source674(spike_out_source[674]),        .spike_out_source675(spike_out_source[675]),        .spike_out_source676(spike_out_source[676]),        .spike_out_source677(spike_out_source[677]),        .spike_out_source678(spike_out_source[678]),        .spike_out_source679(spike_out_source[679]),        .spike_out_source680(spike_out_source[680]),        .spike_out_source681(spike_out_source[681]),        .spike_out_source682(spike_out_source[682]),        .spike_out_source683(spike_out_source[683]),        .spike_out_source684(spike_out_source[684]),        .spike_out_source685(spike_out_source[685]),        .spike_out_source686(spike_out_source[686]),        .spike_out_source687(spike_out_source[687]),        .spike_out_source688(spike_out_source[688]),        .spike_out_source689(spike_out_source[689]),        .spike_out_source690(spike_out_source[690]),        .spike_out_source691(spike_out_source[691]),        .spike_out_source692(spike_out_source[692]),        .spike_out_source693(spike_out_source[693]),        .spike_out_source694(spike_out_source[694]),        .spike_out_source695(spike_out_source[695]),        .spike_out_source696(spike_out_source[696]),        .spike_out_source697(spike_out_source[697]),        .spike_out_source698(spike_out_source[698]),        .spike_out_source699(spike_out_source[699]),        .spike_out_source700(spike_out_source[700]),
        .spike_out_source701(spike_out_source[701]),        .spike_out_source702(spike_out_source[702]),        .spike_out_source703(spike_out_source[703]),        .spike_out_source704(spike_out_source[704]),        .spike_out_source705(spike_out_source[705]),        .spike_out_source706(spike_out_source[706]),        .spike_out_source707(spike_out_source[707]),        .spike_out_source708(spike_out_source[708]),        .spike_out_source709(spike_out_source[709]),        .spike_out_source710(spike_out_source[710]),        .spike_out_source711(spike_out_source[711]),        .spike_out_source712(spike_out_source[712]),        .spike_out_source713(spike_out_source[713]),        .spike_out_source714(spike_out_source[714]),        .spike_out_source715(spike_out_source[715]),        .spike_out_source716(spike_out_source[716]),        .spike_out_source717(spike_out_source[717]),        .spike_out_source718(spike_out_source[718]),        .spike_out_source719(spike_out_source[719]),        .spike_out_source720(spike_out_source[720]),        .spike_out_source721(spike_out_source[721]),        .spike_out_source722(spike_out_source[722]),        .spike_out_source723(spike_out_source[723]),        .spike_out_source724(spike_out_source[724]),        .spike_out_source725(spike_out_source[725]),        .spike_out_source726(spike_out_source[726]),        .spike_out_source727(spike_out_source[727]),        .spike_out_source728(spike_out_source[728]),        .spike_out_source729(spike_out_source[729]),        .spike_out_source730(spike_out_source[730]),        .spike_out_source731(spike_out_source[731]),        .spike_out_source732(spike_out_source[732]),        .spike_out_source733(spike_out_source[733]),        .spike_out_source734(spike_out_source[734]),        .spike_out_source735(spike_out_source[735]),        .spike_out_source736(spike_out_source[736]),        .spike_out_source737(spike_out_source[737]),        .spike_out_source738(spike_out_source[738]),        .spike_out_source739(spike_out_source[739]),        .spike_out_source740(spike_out_source[740]),        .spike_out_source741(spike_out_source[741]),        .spike_out_source742(spike_out_source[742]),        .spike_out_source743(spike_out_source[743]),        .spike_out_source744(spike_out_source[744]),        .spike_out_source745(spike_out_source[745]),        .spike_out_source746(spike_out_source[746]),        .spike_out_source747(spike_out_source[747]),        .spike_out_source748(spike_out_source[748]),        .spike_out_source749(spike_out_source[749]),        .spike_out_source750(spike_out_source[750]),        .spike_out_source751(spike_out_source[751]),        .spike_out_source752(spike_out_source[752]),        .spike_out_source753(spike_out_source[753]),        .spike_out_source754(spike_out_source[754]),        .spike_out_source755(spike_out_source[755]),        .spike_out_source756(spike_out_source[756]),        .spike_out_source757(spike_out_source[757]),        .spike_out_source758(spike_out_source[758]),        .spike_out_source759(spike_out_source[759]),        .spike_out_source760(spike_out_source[760]),        .spike_out_source761(spike_out_source[761]),        .spike_out_source762(spike_out_source[762]),        .spike_out_source763(spike_out_source[763]),        .spike_out_source764(spike_out_source[764]),        .spike_out_source765(spike_out_source[765]),        .spike_out_source766(spike_out_source[766]),        .spike_out_source767(spike_out_source[767]),        .spike_out_source768(spike_out_source[768]),        .spike_out_source769(spike_out_source[769]),        .spike_out_source770(spike_out_source[770]),        .spike_out_source771(spike_out_source[771]),        .spike_out_source772(spike_out_source[772]),        .spike_out_source773(spike_out_source[773]),        .spike_out_source774(spike_out_source[774]),        .spike_out_source775(spike_out_source[775]),        .spike_out_source776(spike_out_source[776]),        .spike_out_source777(spike_out_source[777]),        .spike_out_source778(spike_out_source[778]),        .spike_out_source779(spike_out_source[779]),        .spike_out_source780(spike_out_source[780]),        .spike_out_source781(spike_out_source[781]),        .spike_out_source782(spike_out_source[782]),        .spike_out_source783(spike_out_source[783]),        .spike_out_source784(spike_out_source[784]),        .spike_out_source785(spike_out_source[785]),        .spike_out_source786(spike_out_source[786]),        .spike_out_source787(spike_out_source[787]),        .spike_out_source788(spike_out_source[788]),        .spike_out_source789(spike_out_source[789]),        .spike_out_source790(spike_out_source[790]),        .spike_out_source791(spike_out_source[791]),        .spike_out_source792(spike_out_source[792]),        .spike_out_source793(spike_out_source[793]),        .spike_out_source794(spike_out_source[794]),        .spike_out_source795(spike_out_source[795]),        .spike_out_source796(spike_out_source[796]),        .spike_out_source797(spike_out_source[797]),        .spike_out_source798(spike_out_source[798]),        .spike_out_source799(spike_out_source[799]),        .spike_out_source800(spike_out_source[800]),
        .spike_out_source801(spike_out_source[801]),        .spike_out_source802(spike_out_source[802]),        .spike_out_source803(spike_out_source[803]),        .spike_out_source804(spike_out_source[804]),        .spike_out_source805(spike_out_source[805]),        .spike_out_source806(spike_out_source[806]),        .spike_out_source807(spike_out_source[807]),        .spike_out_source808(spike_out_source[808]),        .spike_out_source809(spike_out_source[809]),        .spike_out_source810(spike_out_source[810]),        .spike_out_source811(spike_out_source[811]),        .spike_out_source812(spike_out_source[812]),        .spike_out_source813(spike_out_source[813]),        .spike_out_source814(spike_out_source[814]),        .spike_out_source815(spike_out_source[815]),        .spike_out_source816(spike_out_source[816]),        .spike_out_source817(spike_out_source[817]),        .spike_out_source818(spike_out_source[818]),        .spike_out_source819(spike_out_source[819]),        .spike_out_source820(spike_out_source[820]),        .spike_out_source821(spike_out_source[821]),        .spike_out_source822(spike_out_source[822]),        .spike_out_source823(spike_out_source[823]),        .spike_out_source824(spike_out_source[824]),        .spike_out_source825(spike_out_source[825]),        .spike_out_source826(spike_out_source[826]),        .spike_out_source827(spike_out_source[827]),        .spike_out_source828(spike_out_source[828]),        .spike_out_source829(spike_out_source[829]),        .spike_out_source830(spike_out_source[830]),        .spike_out_source831(spike_out_source[831]),        .spike_out_source832(spike_out_source[832]),        .spike_out_source833(spike_out_source[833]),        .spike_out_source834(spike_out_source[834]),        .spike_out_source835(spike_out_source[835]),        .spike_out_source836(spike_out_source[836]),        .spike_out_source837(spike_out_source[837]),        .spike_out_source838(spike_out_source[838]),        .spike_out_source839(spike_out_source[839]),        .spike_out_source840(spike_out_source[840]),        .spike_out_source841(spike_out_source[841]),        .spike_out_source842(spike_out_source[842]),        .spike_out_source843(spike_out_source[843]),        .spike_out_source844(spike_out_source[844]),        .spike_out_source845(spike_out_source[845]),        .spike_out_source846(spike_out_source[846]),        .spike_out_source847(spike_out_source[847]),        .spike_out_source848(spike_out_source[848]),        .spike_out_source849(spike_out_source[849]),        .spike_out_source850(spike_out_source[850]),        .spike_out_source851(spike_out_source[851]),        .spike_out_source852(spike_out_source[852]),        .spike_out_source853(spike_out_source[853]),        .spike_out_source854(spike_out_source[854]),        .spike_out_source855(spike_out_source[855]),        .spike_out_source856(spike_out_source[856]),        .spike_out_source857(spike_out_source[857]),        .spike_out_source858(spike_out_source[858]),        .spike_out_source859(spike_out_source[859]),        .spike_out_source860(spike_out_source[860]),        .spike_out_source861(spike_out_source[861]),        .spike_out_source862(spike_out_source[862]),        .spike_out_source863(spike_out_source[863]),        .spike_out_source864(spike_out_source[864]),        .spike_out_source865(spike_out_source[865]),        .spike_out_source866(spike_out_source[866]),        .spike_out_source867(spike_out_source[867]),        .spike_out_source868(spike_out_source[868]),        .spike_out_source869(spike_out_source[869]),        .spike_out_source870(spike_out_source[870]),        .spike_out_source871(spike_out_source[871]),        .spike_out_source872(spike_out_source[872]),        .spike_out_source873(spike_out_source[873]),        .spike_out_source874(spike_out_source[874]),        .spike_out_source875(spike_out_source[875]),        .spike_out_source876(spike_out_source[876]),        .spike_out_source877(spike_out_source[877]),        .spike_out_source878(spike_out_source[878]),        .spike_out_source879(spike_out_source[879]),        .spike_out_source880(spike_out_source[880]),        .spike_out_source881(spike_out_source[881]),        .spike_out_source882(spike_out_source[882]),        .spike_out_source883(spike_out_source[883]),        .spike_out_source884(spike_out_source[884]),        .spike_out_source885(spike_out_source[885]),        .spike_out_source886(spike_out_source[886]),        .spike_out_source887(spike_out_source[887]),        .spike_out_source888(spike_out_source[888]),        .spike_out_source889(spike_out_source[889]),        .spike_out_source890(spike_out_source[890]),        .spike_out_source891(spike_out_source[891]),        .spike_out_source892(spike_out_source[892]),        .spike_out_source893(spike_out_source[893]),        .spike_out_source894(spike_out_source[894]),        .spike_out_source895(spike_out_source[895]),        .spike_out_source896(spike_out_source[896]),        .spike_out_source897(spike_out_source[897]),        .spike_out_source898(spike_out_source[898]),        .spike_out_source899(spike_out_source[899]),        .spike_out_source900(spike_out_source[900]),
        .spike_out_source901(spike_out_source[901]),        .spike_out_source902(spike_out_source[902]),        .spike_out_source903(spike_out_source[903]),        .spike_out_source904(spike_out_source[904]),        .spike_out_source905(spike_out_source[905]),        .spike_out_source906(spike_out_source[906]),        .spike_out_source907(spike_out_source[907]),        .spike_out_source908(spike_out_source[908]),        .spike_out_source909(spike_out_source[909]),        .spike_out_source910(spike_out_source[910]),        .spike_out_source911(spike_out_source[911]),        .spike_out_source912(spike_out_source[912]),        .spike_out_source913(spike_out_source[913]),        .spike_out_source914(spike_out_source[914]),        .spike_out_source915(spike_out_source[915]),        .spike_out_source916(spike_out_source[916]),        .spike_out_source917(spike_out_source[917]),        .spike_out_source918(spike_out_source[918]),        .spike_out_source919(spike_out_source[919]),        .spike_out_source920(spike_out_source[920]),        .spike_out_source921(spike_out_source[921]),        .spike_out_source922(spike_out_source[922]),        .spike_out_source923(spike_out_source[923]),        .spike_out_source924(spike_out_source[924]),        .spike_out_source925(spike_out_source[925]),        .spike_out_source926(spike_out_source[926]),        .spike_out_source927(spike_out_source[927]),        .spike_out_source928(spike_out_source[928]),        .spike_out_source929(spike_out_source[929]),        .spike_out_source930(spike_out_source[930]),        .spike_out_source931(spike_out_source[931]),        .spike_out_source932(spike_out_source[932]),        .spike_out_source933(spike_out_source[933]),        .spike_out_source934(spike_out_source[934]),        .spike_out_source935(spike_out_source[935]),        .spike_out_source936(spike_out_source[936]),        .spike_out_source937(spike_out_source[937]),        .spike_out_source938(spike_out_source[938]),        .spike_out_source939(spike_out_source[939]),        .spike_out_source940(spike_out_source[940]),        .spike_out_source941(spike_out_source[941]),        .spike_out_source942(spike_out_source[942]),        .spike_out_source943(spike_out_source[943]),        .spike_out_source944(spike_out_source[944]),        .spike_out_source945(spike_out_source[945]),        .spike_out_source946(spike_out_source[946]),        .spike_out_source947(spike_out_source[947]),        .spike_out_source948(spike_out_source[948]),        .spike_out_source949(spike_out_source[949]),        .spike_out_source950(spike_out_source[950]),        .spike_out_source951(spike_out_source[951]),        .spike_out_source952(spike_out_source[952]),        .spike_out_source953(spike_out_source[953]),        .spike_out_source954(spike_out_source[954]),        .spike_out_source955(spike_out_source[955]),        .spike_out_source956(spike_out_source[956]),        .spike_out_source957(spike_out_source[957]),        .spike_out_source958(spike_out_source[958]),        .spike_out_source959(spike_out_source[959]),        .spike_out_source960(spike_out_source[960]),        .spike_out_source961(spike_out_source[961]),        .spike_out_source962(spike_out_source[962]),        .spike_out_source963(spike_out_source[963]),        .spike_out_source964(spike_out_source[964]),        .spike_out_source965(spike_out_source[965]),        .spike_out_source966(spike_out_source[966]),        .spike_out_source967(spike_out_source[967]),        .spike_out_source968(spike_out_source[968]),        .spike_out_source969(spike_out_source[969]),        .spike_out_source970(spike_out_source[970]),        .spike_out_source971(spike_out_source[971]),        .spike_out_source972(spike_out_source[972]),        .spike_out_source973(spike_out_source[973]),        .spike_out_source974(spike_out_source[974]),        .spike_out_source975(spike_out_source[975]),        .spike_out_source976(spike_out_source[976]),        .spike_out_source977(spike_out_source[977]),        .spike_out_source978(spike_out_source[978]),        .spike_out_source979(spike_out_source[979]),        .spike_out_source980(spike_out_source[980]),        .spike_out_source981(spike_out_source[981]),        .spike_out_source982(spike_out_source[982]),        .spike_out_source983(spike_out_source[983]),        .spike_out_source984(spike_out_source[984]),        .spike_out_source985(spike_out_source[985]),        .spike_out_source986(spike_out_source[986]),        .spike_out_source987(spike_out_source[987]),        .spike_out_source988(spike_out_source[988]),        .spike_out_source989(spike_out_source[989]),        .spike_out_source990(spike_out_source[990]),        .spike_out_source991(spike_out_source[991]),        .spike_out_source992(spike_out_source[992]),        .spike_out_source993(spike_out_source[993]),        .spike_out_source994(spike_out_source[994]),        .spike_out_source995(spike_out_source[995]),        .spike_out_source996(spike_out_source[996]),        .spike_out_source997(spike_out_source[997]),        .spike_out_source998(spike_out_source[998]),        .spike_out_source999(spike_out_source[999]),        .spike_out_source1000(spike_out_source[1000]),
        .spike_out_source1001(spike_out_source[1001]),        .spike_out_source1002(spike_out_source[1002]),        .spike_out_source1003(spike_out_source[1003]),        .spike_out_source1004(spike_out_source[1004]),        .spike_out_source1005(spike_out_source[1005]),        .spike_out_source1006(spike_out_source[1006]),        .spike_out_source1007(spike_out_source[1007]),        .spike_out_source1008(spike_out_source[1008]),        .spike_out_source1009(spike_out_source[1009]),        .spike_out_source1010(spike_out_source[1010]),        .spike_out_source1011(spike_out_source[1011]),        .spike_out_source1012(spike_out_source[1012]),        .spike_out_source1013(spike_out_source[1013]),        .spike_out_source1014(spike_out_source[1014]),        .spike_out_source1015(spike_out_source[1015]),        .spike_out_source1016(spike_out_source[1016]),        .spike_out_source1017(spike_out_source[1017]),        .spike_out_source1018(spike_out_source[1018]),        .spike_out_source1019(spike_out_source[1019]),        .spike_out_source1020(spike_out_source[1020]),        .spike_out_source1021(spike_out_source[1021]),        .spike_out_source1022(spike_out_source[1022]),        .spike_out_source1023(spike_out_source[1023])
endmodule
