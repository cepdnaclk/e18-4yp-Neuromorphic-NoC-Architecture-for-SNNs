`timescale 1ns/100ps
// `include "potential_decay.v"
// `include "mac.v"
// `include "Addition_Subtraction.v"
// `include "potential_adder.v"
// `include "network_interface.v"
// `include "Multiplication.v"

module testbench;

    parameter number_of_units = 1024;
    parameter number_of_neurons=10;                         //initiailize number of neurons
    reg CLK;                                                //clock
    reg clear;                                              //clear to start timestep
    reg[3:0] decay_rate;                                    //define decay rate
    reg[3:0] CLK_count;                                     //counter for clocks

    reg[11:0] source_addresses[0:number_of_units-1];          //write her simulate spike packets by sending source addresses
    reg[159:0] weights_arrays[0:number_of_units-1];           //initialize store weights of the connections
    reg[59:0] source_addresses_arrays[0:number_of_units-1];   //initialize connection by writing source addresses to the accumulators
                                                              //12 bits * 5 max connections
    reg[11:0] neuron_addresses[0:number_of_units-1];          //initialize with neuron addresses
    reg[31:0] membrane_potential[0:number_of_units-1];        //initialize membrane potential values
    reg[31:0] v_threshold[0:number_of_units-1];               //threshold values
    reg[359:0] downstream_connections_initialization;           //input to initialize the dowanstream connections
                                                                //12bits * 10 SNN neurons * 3 connections per nueron
                                                                
    reg[119:0] neuron_addresses_initialization;                 //input to initialize the neruon addresses
                                                                //12 bits * 10 SNN neurons
    reg[54:0] connection_pointer_initialization;                //input to initialize the connection pointers
                                                                //11 row pointer elements * 5 bits (to represent 30 connections)
    reg[11:0] spike_origin;                                     //to store the nueron address from the arrived packet
    reg[11:0] spike_destination;                                //to store source address from the arrived packet
    
    reg[1:0] model;
    reg[31:0]a, b, c, d, u_initialize;      //for izhikevich model
    
    wire[31:0] results_mac[0:number_of_units-1];                 //store results from the mac
    wire[31:0] results_potential_decay[0:number_of_units-1];     //store results of potential decay
    wire[31:0] final_potential[0:number_of_units-1];             //potential form the potential adder
    wire spike[0:number_of_units-1];                              //spike signifier from potential decay
    // wire[23:0] packet1, packet2, packet3, packet4, packet5, packet6, packet7, packet8, packet9,
    //         packet10, packet11, packet12, packet13, packet14, packet15, packet16, packet17, packet18,
    //         packet19, packet20, packet21;                          //packet containing neuron address and sources address

    //intermediate wires to hold the output of the network interface
    wire[11:0] spike_out_source[0:number_of_units-1];
    
    // wires and registers needed for the fifo buffers
    reg rst_n;
    reg wr_en;
    reg rd_en;
    wire [11:0] rd_data [1023:0];
    wire empty [1023:0];
    wire full [1023:0];

    // create 1024 FIFO buffers
    // between the network interface and mac
    genvar i;
    generate
        for (i = 0; i < number_of_units; i = i+1) begin
            async_fifo_copy fifo1 (
                .rd_clk(clear),
                .rst_n(rst_n),
                // .wr_en(~clear),
                .wr_en(wr_en),
                .wr_data(spike_out_source[i]),      // send the input from ni to the fifo
                .rd_en(clear),
                .rd_data(rd_data[i]),               // send the read source addresses to the mac
                .empty(empty[i]),
                .full(full[i])
            );
        end
    endgenerate
    


    //generate 1024 potential decay units
    generate
        for(i=0; i<number_of_units; i=i+1) begin
            potential_decay pd(
                .CLK(CLK),
                .clear(clear),
                .model(model),
                .neuron_address_initialization(neuron_addresses[i]),
                .decay_rate(decay_rate),
                .membrane_potential_initialization(membrane_potential[i]),
                .output_potential_decay(results_potential_decay[i]),
                .new_potential(final_potential[i])
            );
        end
    endgenerate

    //generate 1024 accumulators
    generate
        for(i=0; i<number_of_units; i=i+1) begin
            mac m(
                .CLK(CLK),
                .neuron_address(neuron_addresses[i]),
                // .source_address(spike_out_source[i]),
                .source_address(rd_data[i]),
                .weights_array(weights_arrays[i]),
                .source_addresses_array(source_addresses_arrays[i]),
                .clear(clear),
                .mult_output(results_mac[i])
            );
        end
    endgenerate

    //genrate corresponding 1024 potential adders
    generate
        for(i=0; i<number_of_units; i=i+1) begin
            potential_adder pa(
                .clear(clear),
                .v_threshold(v_threshold[i]),
                .input_weight(results_mac[i]),
                .decayed_potential(results_potential_decay[i]),
                .model(model),
                .a(a),
                .b(b),
                .c(c),
                .d(d),
                .u_initialize(u_initialize),
                .final_potential(final_potential[i]),
                .spike(spike[i])
            );
        end
    endgenerate

    //network interface initialisation
    network_interface_new ni1(
        .CLK(CLK),
        .clear(clear),
        .spike0(spike[0]),
        .spike1(spike[1]),        .spike2(spike[2]),        .spike3(spike[3]),        .spike4(spike[4]),        .spike5(spike[5]),        .spike6(spike[6]),        .spike7(spike[7]),        .spike8(spike[8]),        .spike9(spike[9]),        .spike10(spike[10]),        .spike11(spike[11]),        .spike12(spike[12]),        .spike13(spike[13]),        .spike14(spike[14]),        .spike15(spike[15]),        .spike16(spike[16]),        .spike17(spike[17]),        .spike18(spike[18]),        .spike19(spike[19]),        .spike20(spike[20]),        .spike21(spike[21]),        .spike22(spike[22]),        .spike23(spike[23]),        .spike24(spike[24]),        .spike25(spike[25]),        .spike26(spike[26]),        .spike27(spike[27]),        .spike28(spike[28]),        .spike29(spike[29]),        .spike30(spike[30]),        .spike31(spike[31]),        .spike32(spike[32]),        .spike33(spike[33]),        .spike34(spike[34]),        .spike35(spike[35]),        .spike36(spike[36]),        .spike37(spike[37]),        .spike38(spike[38]),        .spike39(spike[39]),        .spike40(spike[40]),        .spike41(spike[41]),        .spike42(spike[42]),        .spike43(spike[43]),        .spike44(spike[44]),        .spike45(spike[45]),        .spike46(spike[46]),        .spike47(spike[47]),        .spike48(spike[48]),        .spike49(spike[49]),        .spike50(spike[50]),        .spike51(spike[51]),        .spike52(spike[52]),        .spike53(spike[53]),        .spike54(spike[54]),        .spike55(spike[55]),        .spike56(spike[56]),        .spike57(spike[57]),        .spike58(spike[58]),        .spike59(spike[59]),        .spike60(spike[60]),        .spike61(spike[61]),        .spike62(spike[62]),        .spike63(spike[63]),        .spike64(spike[64]),        .spike65(spike[65]),        .spike66(spike[66]),        .spike67(spike[67]),        .spike68(spike[68]),        .spike69(spike[69]),        .spike70(spike[70]),        .spike71(spike[71]),        .spike72(spike[72]),        .spike73(spike[73]),        .spike74(spike[74]),        .spike75(spike[75]),        .spike76(spike[76]),        .spike77(spike[77]),        .spike78(spike[78]),        .spike79(spike[79]),        .spike80(spike[80]),        .spike81(spike[81]),        .spike82(spike[82]),        .spike83(spike[83]),        .spike84(spike[84]),        .spike85(spike[85]),        .spike86(spike[86]),        .spike87(spike[87]),        .spike88(spike[88]),        .spike89(spike[89]),        .spike90(spike[90]),        .spike91(spike[91]),        .spike92(spike[92]),        .spike93(spike[93]),        .spike94(spike[94]),        .spike95(spike[95]),        .spike96(spike[96]),        .spike97(spike[97]),        .spike98(spike[98]),        .spike99(spike[99]),        .spike100(spike[100]),
        .spike101(spike[101]),        .spike102(spike[102]),        .spike103(spike[103]),        .spike104(spike[104]),        .spike105(spike[105]),        .spike106(spike[106]),        .spike107(spike[107]),        .spike108(spike[108]),        .spike109(spike[109]),        .spike110(spike[110]),        .spike111(spike[111]),        .spike112(spike[112]),        .spike113(spike[113]),        .spike114(spike[114]),        .spike115(spike[115]),        .spike116(spike[116]),        .spike117(spike[117]),        .spike118(spike[118]),        .spike119(spike[119]),        .spike120(spike[120]),        .spike121(spike[121]),        .spike122(spike[122]),        .spike123(spike[123]),        .spike124(spike[124]),        .spike125(spike[125]),        .spike126(spike[126]),        .spike127(spike[127]),        .spike128(spike[128]),        .spike129(spike[129]),        .spike130(spike[130]),        .spike131(spike[131]),        .spike132(spike[132]),        .spike133(spike[133]),        .spike134(spike[134]),        .spike135(spike[135]),        .spike136(spike[136]),        .spike137(spike[137]),        .spike138(spike[138]),        .spike139(spike[139]),        .spike140(spike[140]),        .spike141(spike[141]),        .spike142(spike[142]),        .spike143(spike[143]),        .spike144(spike[144]),        .spike145(spike[145]),        .spike146(spike[146]),        .spike147(spike[147]),        .spike148(spike[148]),        .spike149(spike[149]),        .spike150(spike[150]),        .spike151(spike[151]),        .spike152(spike[152]),        .spike153(spike[153]),        .spike154(spike[154]),        .spike155(spike[155]),        .spike156(spike[156]),        .spike157(spike[157]),        .spike158(spike[158]),        .spike159(spike[159]),        .spike160(spike[160]),        .spike161(spike[161]),        .spike162(spike[162]),        .spike163(spike[163]),        .spike164(spike[164]),        .spike165(spike[165]),        .spike166(spike[166]),        .spike167(spike[167]),        .spike168(spike[168]),        .spike169(spike[169]),        .spike170(spike[170]),        .spike171(spike[171]),        .spike172(spike[172]),        .spike173(spike[173]),        .spike174(spike[174]),        .spike175(spike[175]),        .spike176(spike[176]),        .spike177(spike[177]),        .spike178(spike[178]),        .spike179(spike[179]),        .spike180(spike[180]),        .spike181(spike[181]),        .spike182(spike[182]),        .spike183(spike[183]),        .spike184(spike[184]),        .spike185(spike[185]),        .spike186(spike[186]),        .spike187(spike[187]),        .spike188(spike[188]),        .spike189(spike[189]),        .spike190(spike[190]),        .spike191(spike[191]),        .spike192(spike[192]),        .spike193(spike[193]),        .spike194(spike[194]),        .spike195(spike[195]),        .spike196(spike[196]),        .spike197(spike[197]),        .spike198(spike[198]),        .spike199(spike[199]),        .spike200(spike[200]),
        .spike201(spike[201]),        .spike202(spike[202]),        .spike203(spike[203]),        .spike204(spike[204]),        .spike205(spike[205]),        .spike206(spike[206]),        .spike207(spike[207]),        .spike208(spike[208]),        .spike209(spike[209]),        .spike210(spike[210]),        .spike211(spike[211]),        .spike212(spike[212]),        .spike213(spike[213]),        .spike214(spike[214]),        .spike215(spike[215]),        .spike216(spike[216]),        .spike217(spike[217]),        .spike218(spike[218]),        .spike219(spike[219]),        .spike220(spike[220]),        .spike221(spike[221]),        .spike222(spike[222]),        .spike223(spike[223]),        .spike224(spike[224]),        .spike225(spike[225]),        .spike226(spike[226]),        .spike227(spike[227]),        .spike228(spike[228]),        .spike229(spike[229]),        .spike230(spike[230]),        .spike231(spike[231]),        .spike232(spike[232]),        .spike233(spike[233]),        .spike234(spike[234]),        .spike235(spike[235]),        .spike236(spike[236]),        .spike237(spike[237]),        .spike238(spike[238]),        .spike239(spike[239]),        .spike240(spike[240]),        .spike241(spike[241]),        .spike242(spike[242]),        .spike243(spike[243]),        .spike244(spike[244]),        .spike245(spike[245]),        .spike246(spike[246]),        .spike247(spike[247]),        .spike248(spike[248]),        .spike249(spike[249]),        .spike250(spike[250]),        .spike251(spike[251]),        .spike252(spike[252]),        .spike253(spike[253]),        .spike254(spike[254]),        .spike255(spike[255]),        .spike256(spike[256]),        .spike257(spike[257]),        .spike258(spike[258]),        .spike259(spike[259]),        .spike260(spike[260]),        .spike261(spike[261]),        .spike262(spike[262]),        .spike263(spike[263]),        .spike264(spike[264]),        .spike265(spike[265]),        .spike266(spike[266]),        .spike267(spike[267]),        .spike268(spike[268]),        .spike269(spike[269]),        .spike270(spike[270]),        .spike271(spike[271]),        .spike272(spike[272]),        .spike273(spike[273]),        .spike274(spike[274]),        .spike275(spike[275]),        .spike276(spike[276]),        .spike277(spike[277]),        .spike278(spike[278]),        .spike279(spike[279]),        .spike280(spike[280]),        .spike281(spike[281]),        .spike282(spike[282]),        .spike283(spike[283]),        .spike284(spike[284]),        .spike285(spike[285]),        .spike286(spike[286]),        .spike287(spike[287]),        .spike288(spike[288]),        .spike289(spike[289]),        .spike290(spike[290]),        .spike291(spike[291]),        .spike292(spike[292]),        .spike293(spike[293]),        .spike294(spike[294]),        .spike295(spike[295]),        .spike296(spike[296]),        .spike297(spike[297]),        .spike298(spike[298]),        .spike299(spike[299]),        .spike300(spike[300]),
        .spike301(spike[301]),        .spike302(spike[302]),        .spike303(spike[303]),        .spike304(spike[304]),        .spike305(spike[305]),        .spike306(spike[306]),        .spike307(spike[307]),        .spike308(spike[308]),        .spike309(spike[309]),        .spike310(spike[310]),        .spike311(spike[311]),        .spike312(spike[312]),        .spike313(spike[313]),        .spike314(spike[314]),        .spike315(spike[315]),        .spike316(spike[316]),        .spike317(spike[317]),        .spike318(spike[318]),        .spike319(spike[319]),        .spike320(spike[320]),        .spike321(spike[321]),        .spike322(spike[322]),        .spike323(spike[323]),        .spike324(spike[324]),        .spike325(spike[325]),        .spike326(spike[326]),        .spike327(spike[327]),        .spike328(spike[328]),        .spike329(spike[329]),        .spike330(spike[330]),        .spike331(spike[331]),        .spike332(spike[332]),        .spike333(spike[333]),        .spike334(spike[334]),        .spike335(spike[335]),        .spike336(spike[336]),        .spike337(spike[337]),        .spike338(spike[338]),        .spike339(spike[339]),        .spike340(spike[340]),        .spike341(spike[341]),        .spike342(spike[342]),        .spike343(spike[343]),        .spike344(spike[344]),        .spike345(spike[345]),        .spike346(spike[346]),        .spike347(spike[347]),        .spike348(spike[348]),        .spike349(spike[349]),        .spike350(spike[350]),        .spike351(spike[351]),        .spike352(spike[352]),        .spike353(spike[353]),        .spike354(spike[354]),        .spike355(spike[355]),        .spike356(spike[356]),        .spike357(spike[357]),        .spike358(spike[358]),        .spike359(spike[359]),        .spike360(spike[360]),        .spike361(spike[361]),        .spike362(spike[362]),        .spike363(spike[363]),        .spike364(spike[364]),        .spike365(spike[365]),        .spike366(spike[366]),        .spike367(spike[367]),        .spike368(spike[368]),        .spike369(spike[369]),        .spike370(spike[370]),        .spike371(spike[371]),        .spike372(spike[372]),        .spike373(spike[373]),        .spike374(spike[374]),        .spike375(spike[375]),        .spike376(spike[376]),        .spike377(spike[377]),        .spike378(spike[378]),        .spike379(spike[379]),        .spike380(spike[380]),        .spike381(spike[381]),        .spike382(spike[382]),        .spike383(spike[383]),        .spike384(spike[384]),        .spike385(spike[385]),        .spike386(spike[386]),        .spike387(spike[387]),        .spike388(spike[388]),        .spike389(spike[389]),        .spike390(spike[390]),        .spike391(spike[391]),        .spike392(spike[392]),        .spike393(spike[393]),        .spike394(spike[394]),        .spike395(spike[395]),        .spike396(spike[396]),        .spike397(spike[397]),        .spike398(spike[398]),        .spike399(spike[399]),        .spike400(spike[400]),
        .spike401(spike[401]),        .spike402(spike[402]),        .spike403(spike[403]),        .spike404(spike[404]),        .spike405(spike[405]),        .spike406(spike[406]),        .spike407(spike[407]),        .spike408(spike[408]),        .spike409(spike[409]),        .spike410(spike[410]),        .spike411(spike[411]),        .spike412(spike[412]),        .spike413(spike[413]),        .spike414(spike[414]),        .spike415(spike[415]),        .spike416(spike[416]),        .spike417(spike[417]),        .spike418(spike[418]),        .spike419(spike[419]),        .spike420(spike[420]),        .spike421(spike[421]),        .spike422(spike[422]),        .spike423(spike[423]),        .spike424(spike[424]),        .spike425(spike[425]),        .spike426(spike[426]),        .spike427(spike[427]),        .spike428(spike[428]),        .spike429(spike[429]),        .spike430(spike[430]),        .spike431(spike[431]),        .spike432(spike[432]),        .spike433(spike[433]),        .spike434(spike[434]),        .spike435(spike[435]),        .spike436(spike[436]),        .spike437(spike[437]),        .spike438(spike[438]),        .spike439(spike[439]),        .spike440(spike[440]),        .spike441(spike[441]),        .spike442(spike[442]),        .spike443(spike[443]),        .spike444(spike[444]),        .spike445(spike[445]),        .spike446(spike[446]),        .spike447(spike[447]),        .spike448(spike[448]),        .spike449(spike[449]),        .spike450(spike[450]),        .spike451(spike[451]),        .spike452(spike[452]),        .spike453(spike[453]),        .spike454(spike[454]),        .spike455(spike[455]),        .spike456(spike[456]),        .spike457(spike[457]),        .spike458(spike[458]),        .spike459(spike[459]),        .spike460(spike[460]),        .spike461(spike[461]),        .spike462(spike[462]),        .spike463(spike[463]),        .spike464(spike[464]),        .spike465(spike[465]),        .spike466(spike[466]),        .spike467(spike[467]),        .spike468(spike[468]),        .spike469(spike[469]),        .spike470(spike[470]),        .spike471(spike[471]),        .spike472(spike[472]),        .spike473(spike[473]),        .spike474(spike[474]),        .spike475(spike[475]),        .spike476(spike[476]),        .spike477(spike[477]),        .spike478(spike[478]),        .spike479(spike[479]),        .spike480(spike[480]),        .spike481(spike[481]),        .spike482(spike[482]),        .spike483(spike[483]),        .spike484(spike[484]),        .spike485(spike[485]),        .spike486(spike[486]),        .spike487(spike[487]),        .spike488(spike[488]),        .spike489(spike[489]),        .spike490(spike[490]),        .spike491(spike[491]),        .spike492(spike[492]),        .spike493(spike[493]),        .spike494(spike[494]),        .spike495(spike[495]),        .spike496(spike[496]),        .spike497(spike[497]),        .spike498(spike[498]),        .spike499(spike[499]),        .spike500(spike[500]),
        .spike501(spike[501]),        .spike502(spike[502]),        .spike503(spike[503]),        .spike504(spike[504]),        .spike505(spike[505]),        .spike506(spike[506]),        .spike507(spike[507]),        .spike508(spike[508]),        .spike509(spike[509]),        .spike510(spike[510]),        .spike511(spike[511]),        .spike512(spike[512]),        .spike513(spike[513]),        .spike514(spike[514]),        .spike515(spike[515]),        .spike516(spike[516]),        .spike517(spike[517]),        .spike518(spike[518]),        .spike519(spike[519]),        .spike520(spike[520]),        .spike521(spike[521]),        .spike522(spike[522]),        .spike523(spike[523]),        .spike524(spike[524]),        .spike525(spike[525]),        .spike526(spike[526]),        .spike527(spike[527]),        .spike528(spike[528]),        .spike529(spike[529]),        .spike530(spike[530]),        .spike531(spike[531]),        .spike532(spike[532]),        .spike533(spike[533]),        .spike534(spike[534]),        .spike535(spike[535]),        .spike536(spike[536]),        .spike537(spike[537]),        .spike538(spike[538]),        .spike539(spike[539]),        .spike540(spike[540]),        .spike541(spike[541]),        .spike542(spike[542]),        .spike543(spike[543]),        .spike544(spike[544]),        .spike545(spike[545]),        .spike546(spike[546]),        .spike547(spike[547]),        .spike548(spike[548]),        .spike549(spike[549]),        .spike550(spike[550]),        .spike551(spike[551]),        .spike552(spike[552]),        .spike553(spike[553]),        .spike554(spike[554]),        .spike555(spike[555]),        .spike556(spike[556]),        .spike557(spike[557]),        .spike558(spike[558]),        .spike559(spike[559]),        .spike560(spike[560]),        .spike561(spike[561]),        .spike562(spike[562]),        .spike563(spike[563]),        .spike564(spike[564]),        .spike565(spike[565]),        .spike566(spike[566]),        .spike567(spike[567]),        .spike568(spike[568]),        .spike569(spike[569]),        .spike570(spike[570]),        .spike571(spike[571]),        .spike572(spike[572]),        .spike573(spike[573]),        .spike574(spike[574]),        .spike575(spike[575]),        .spike576(spike[576]),        .spike577(spike[577]),        .spike578(spike[578]),        .spike579(spike[579]),        .spike580(spike[580]),        .spike581(spike[581]),        .spike582(spike[582]),        .spike583(spike[583]),        .spike584(spike[584]),        .spike585(spike[585]),        .spike586(spike[586]),        .spike587(spike[587]),        .spike588(spike[588]),        .spike589(spike[589]),        .spike590(spike[590]),        .spike591(spike[591]),        .spike592(spike[592]),        .spike593(spike[593]),        .spike594(spike[594]),        .spike595(spike[595]),        .spike596(spike[596]),        .spike597(spike[597]),        .spike598(spike[598]),        .spike599(spike[599]),        .spike600(spike[600]),
        .spike601(spike[601]),        .spike602(spike[602]),        .spike603(spike[603]),        .spike604(spike[604]),        .spike605(spike[605]),        .spike606(spike[606]),        .spike607(spike[607]),        .spike608(spike[608]),        .spike609(spike[609]),        .spike610(spike[610]),        .spike611(spike[611]),        .spike612(spike[612]),        .spike613(spike[613]),        .spike614(spike[614]),        .spike615(spike[615]),        .spike616(spike[616]),        .spike617(spike[617]),        .spike618(spike[618]),        .spike619(spike[619]),        .spike620(spike[620]),        .spike621(spike[621]),        .spike622(spike[622]),        .spike623(spike[623]),        .spike624(spike[624]),        .spike625(spike[625]),        .spike626(spike[626]),        .spike627(spike[627]),        .spike628(spike[628]),        .spike629(spike[629]),        .spike630(spike[630]),        .spike631(spike[631]),        .spike632(spike[632]),        .spike633(spike[633]),        .spike634(spike[634]),        .spike635(spike[635]),        .spike636(spike[636]),        .spike637(spike[637]),        .spike638(spike[638]),        .spike639(spike[639]),        .spike640(spike[640]),        .spike641(spike[641]),        .spike642(spike[642]),        .spike643(spike[643]),        .spike644(spike[644]),        .spike645(spike[645]),        .spike646(spike[646]),        .spike647(spike[647]),        .spike648(spike[648]),        .spike649(spike[649]),        .spike650(spike[650]),        .spike651(spike[651]),        .spike652(spike[652]),        .spike653(spike[653]),        .spike654(spike[654]),        .spike655(spike[655]),        .spike656(spike[656]),        .spike657(spike[657]),        .spike658(spike[658]),        .spike659(spike[659]),        .spike660(spike[660]),        .spike661(spike[661]),        .spike662(spike[662]),        .spike663(spike[663]),        .spike664(spike[664]),        .spike665(spike[665]),        .spike666(spike[666]),        .spike667(spike[667]),        .spike668(spike[668]),        .spike669(spike[669]),        .spike670(spike[670]),        .spike671(spike[671]),        .spike672(spike[672]),        .spike673(spike[673]),        .spike674(spike[674]),        .spike675(spike[675]),        .spike676(spike[676]),        .spike677(spike[677]),        .spike678(spike[678]),        .spike679(spike[679]),        .spike680(spike[680]),        .spike681(spike[681]),        .spike682(spike[682]),        .spike683(spike[683]),        .spike684(spike[684]),        .spike685(spike[685]),        .spike686(spike[686]),        .spike687(spike[687]),        .spike688(spike[688]),        .spike689(spike[689]),        .spike690(spike[690]),        .spike691(spike[691]),        .spike692(spike[692]),        .spike693(spike[693]),        .spike694(spike[694]),        .spike695(spike[695]),        .spike696(spike[696]),        .spike697(spike[697]),        .spike698(spike[698]),        .spike699(spike[699]),        .spike700(spike[700]),
        .spike701(spike[701]),        .spike702(spike[702]),        .spike703(spike[703]),        .spike704(spike[704]),        .spike705(spike[705]),        .spike706(spike[706]),        .spike707(spike[707]),        .spike708(spike[708]),        .spike709(spike[709]),        .spike710(spike[710]),        .spike711(spike[711]),        .spike712(spike[712]),        .spike713(spike[713]),        .spike714(spike[714]),        .spike715(spike[715]),        .spike716(spike[716]),        .spike717(spike[717]),        .spike718(spike[718]),        .spike719(spike[719]),        .spike720(spike[720]),        .spike721(spike[721]),        .spike722(spike[722]),        .spike723(spike[723]),        .spike724(spike[724]),        .spike725(spike[725]),        .spike726(spike[726]),        .spike727(spike[727]),        .spike728(spike[728]),        .spike729(spike[729]),        .spike730(spike[730]),        .spike731(spike[731]),        .spike732(spike[732]),        .spike733(spike[733]),        .spike734(spike[734]),        .spike735(spike[735]),        .spike736(spike[736]),        .spike737(spike[737]),        .spike738(spike[738]),        .spike739(spike[739]),        .spike740(spike[740]),        .spike741(spike[741]),        .spike742(spike[742]),        .spike743(spike[743]),        .spike744(spike[744]),        .spike745(spike[745]),        .spike746(spike[746]),        .spike747(spike[747]),        .spike748(spike[748]),        .spike749(spike[749]),        .spike750(spike[750]),        .spike751(spike[751]),        .spike752(spike[752]),        .spike753(spike[753]),        .spike754(spike[754]),        .spike755(spike[755]),        .spike756(spike[756]),        .spike757(spike[757]),        .spike758(spike[758]),        .spike759(spike[759]),        .spike760(spike[760]),        .spike761(spike[761]),        .spike762(spike[762]),        .spike763(spike[763]),        .spike764(spike[764]),        .spike765(spike[765]),        .spike766(spike[766]),        .spike767(spike[767]),        .spike768(spike[768]),        .spike769(spike[769]),        .spike770(spike[770]),        .spike771(spike[771]),        .spike772(spike[772]),        .spike773(spike[773]),        .spike774(spike[774]),        .spike775(spike[775]),        .spike776(spike[776]),        .spike777(spike[777]),        .spike778(spike[778]),        .spike779(spike[779]),        .spike780(spike[780]),        .spike781(spike[781]),        .spike782(spike[782]),        .spike783(spike[783]),        .spike784(spike[784]),        .spike785(spike[785]),        .spike786(spike[786]),        .spike787(spike[787]),        .spike788(spike[788]),        .spike789(spike[789]),        .spike790(spike[790]),        .spike791(spike[791]),        .spike792(spike[792]),        .spike793(spike[793]),        .spike794(spike[794]),        .spike795(spike[795]),        .spike796(spike[796]),        .spike797(spike[797]),        .spike798(spike[798]),        .spike799(spike[799]),        .spike800(spike[800]),
        .spike801(spike[801]),        .spike802(spike[802]),        .spike803(spike[803]),        .spike804(spike[804]),        .spike805(spike[805]),        .spike806(spike[806]),        .spike807(spike[807]),        .spike808(spike[808]),        .spike809(spike[809]),        .spike810(spike[810]),        .spike811(spike[811]),        .spike812(spike[812]),        .spike813(spike[813]),        .spike814(spike[814]),        .spike815(spike[815]),        .spike816(spike[816]),        .spike817(spike[817]),        .spike818(spike[818]),        .spike819(spike[819]),        .spike820(spike[820]),        .spike821(spike[821]),        .spike822(spike[822]),        .spike823(spike[823]),        .spike824(spike[824]),        .spike825(spike[825]),        .spike826(spike[826]),        .spike827(spike[827]),        .spike828(spike[828]),        .spike829(spike[829]),        .spike830(spike[830]),        .spike831(spike[831]),        .spike832(spike[832]),        .spike833(spike[833]),        .spike834(spike[834]),        .spike835(spike[835]),        .spike836(spike[836]),        .spike837(spike[837]),        .spike838(spike[838]),        .spike839(spike[839]),        .spike840(spike[840]),        .spike841(spike[841]),        .spike842(spike[842]),        .spike843(spike[843]),        .spike844(spike[844]),        .spike845(spike[845]),        .spike846(spike[846]),        .spike847(spike[847]),        .spike848(spike[848]),        .spike849(spike[849]),        .spike850(spike[850]),        .spike851(spike[851]),        .spike852(spike[852]),        .spike853(spike[853]),        .spike854(spike[854]),        .spike855(spike[855]),        .spike856(spike[856]),        .spike857(spike[857]),        .spike858(spike[858]),        .spike859(spike[859]),        .spike860(spike[860]),        .spike861(spike[861]),        .spike862(spike[862]),        .spike863(spike[863]),        .spike864(spike[864]),        .spike865(spike[865]),        .spike866(spike[866]),        .spike867(spike[867]),        .spike868(spike[868]),        .spike869(spike[869]),        .spike870(spike[870]),        .spike871(spike[871]),        .spike872(spike[872]),        .spike873(spike[873]),        .spike874(spike[874]),        .spike875(spike[875]),        .spike876(spike[876]),        .spike877(spike[877]),        .spike878(spike[878]),        .spike879(spike[879]),        .spike880(spike[880]),        .spike881(spike[881]),        .spike882(spike[882]),        .spike883(spike[883]),        .spike884(spike[884]),        .spike885(spike[885]),        .spike886(spike[886]),        .spike887(spike[887]),        .spike888(spike[888]),        .spike889(spike[889]),        .spike890(spike[890]),        .spike891(spike[891]),        .spike892(spike[892]),        .spike893(spike[893]),        .spike894(spike[894]),        .spike895(spike[895]),        .spike896(spike[896]),        .spike897(spike[897]),        .spike898(spike[898]),        .spike899(spike[899]),        .spike900(spike[900]),
        .spike901(spike[901]),        .spike902(spike[902]),        .spike903(spike[903]),        .spike904(spike[904]),        .spike905(spike[905]),        .spike906(spike[906]),        .spike907(spike[907]),        .spike908(spike[908]),        .spike909(spike[909]),        .spike910(spike[910]),        .spike911(spike[911]),        .spike912(spike[912]),        .spike913(spike[913]),        .spike914(spike[914]),        .spike915(spike[915]),        .spike916(spike[916]),        .spike917(spike[917]),        .spike918(spike[918]),        .spike919(spike[919]),        .spike920(spike[920]),        .spike921(spike[921]),        .spike922(spike[922]),        .spike923(spike[923]),        .spike924(spike[924]),        .spike925(spike[925]),        .spike926(spike[926]),        .spike927(spike[927]),        .spike928(spike[928]),        .spike929(spike[929]),        .spike930(spike[930]),        .spike931(spike[931]),        .spike932(spike[932]),        .spike933(spike[933]),        .spike934(spike[934]),        .spike935(spike[935]),        .spike936(spike[936]),        .spike937(spike[937]),        .spike938(spike[938]),        .spike939(spike[939]),        .spike940(spike[940]),        .spike941(spike[941]),        .spike942(spike[942]),        .spike943(spike[943]),        .spike944(spike[944]),        .spike945(spike[945]),        .spike946(spike[946]),        .spike947(spike[947]),        .spike948(spike[948]),        .spike949(spike[949]),        .spike950(spike[950]),        .spike951(spike[951]),        .spike952(spike[952]),        .spike953(spike[953]),        .spike954(spike[954]),        .spike955(spike[955]),        .spike956(spike[956]),        .spike957(spike[957]),        .spike958(spike[958]),        .spike959(spike[959]),        .spike960(spike[960]),        .spike961(spike[961]),        .spike962(spike[962]),        .spike963(spike[963]),        .spike964(spike[964]),        .spike965(spike[965]),        .spike966(spike[966]),        .spike967(spike[967]),        .spike968(spike[968]),        .spike969(spike[969]),        .spike970(spike[970]),        .spike971(spike[971]),        .spike972(spike[972]),        .spike973(spike[973]),        .spike974(spike[974]),        .spike975(spike[975]),        .spike976(spike[976]),        .spike977(spike[977]),        .spike978(spike[978]),        .spike979(spike[979]),        .spike980(spike[980]),        .spike981(spike[981]),        .spike982(spike[982]),        .spike983(spike[983]),        .spike984(spike[984]),        .spike985(spike[985]),        .spike986(spike[986]),        .spike987(spike[987]),        .spike988(spike[988]),        .spike989(spike[989]),        .spike990(spike[990]),        .spike991(spike[991]),        .spike992(spike[992]),        .spike993(spike[993]),        .spike994(spike[994]),        .spike995(spike[995]),        .spike996(spike[996]),        .spike997(spike[997]),        .spike998(spike[998]),        .spike999(spike[999]),        .spike1000(spike[1000]),
        .spike1001(spike[1001]),        .spike1002(spike[1002]),        .spike1003(spike[1003]),        .spike1004(spike[1004]),        .spike1005(spike[1005]),        .spike1006(spike[1006]),        .spike1007(spike[1007]),        .spike1008(spike[1008]),        .spike1009(spike[1009]),        .spike1010(spike[1010]),        .spike1011(spike[1011]),        .spike1012(spike[1012]),        .spike1013(spike[1013]),        .spike1014(spike[1014]),        .spike1015(spike[1015]),        .spike1016(spike[1016]),        .spike1017(spike[1017]),        .spike1018(spike[1018]),        .spike1019(spike[1019]),        .spike1020(spike[1020]),        .spike1021(spike[1021]),        .spike1022(spike[1022]),        .spike1023(spike[1023]),
        .neuron_addresses_initialization(neuron_addresses_initialization),
        .connection_pointer_initialization(connection_pointer_initialization),           //input to initialize the connection pointers
        .downstream_connections_initialization(downstream_connections_initialization),    //input to initialize the dowanstream connections
        .spike_out_source0(spike_out_source[0]),            .spike_out_source1(spike_out_source[1]),        .spike_out_source2(spike_out_source[2]),        .spike_out_source3(spike_out_source[3]),        .spike_out_source4(spike_out_source[4]),        .spike_out_source5(spike_out_source[5]),        .spike_out_source6(spike_out_source[6]),        .spike_out_source7(spike_out_source[7]),        .spike_out_source8(spike_out_source[8]),        .spike_out_source9(spike_out_source[9]),        .spike_out_source10(spike_out_source[10]),        .spike_out_source11(spike_out_source[11]),        .spike_out_source12(spike_out_source[12]),        .spike_out_source13(spike_out_source[13]),        .spike_out_source14(spike_out_source[14]),        .spike_out_source15(spike_out_source[15]),        .spike_out_source16(spike_out_source[16]),        .spike_out_source17(spike_out_source[17]),        .spike_out_source18(spike_out_source[18]),        .spike_out_source19(spike_out_source[19]),        .spike_out_source20(spike_out_source[20]),        .spike_out_source21(spike_out_source[21]),        .spike_out_source22(spike_out_source[22]),        .spike_out_source23(spike_out_source[23]),        .spike_out_source24(spike_out_source[24]),        .spike_out_source25(spike_out_source[25]),        .spike_out_source26(spike_out_source[26]),        .spike_out_source27(spike_out_source[27]),        .spike_out_source28(spike_out_source[28]),        .spike_out_source29(spike_out_source[29]),        .spike_out_source30(spike_out_source[30]),        .spike_out_source31(spike_out_source[31]),        .spike_out_source32(spike_out_source[32]),        .spike_out_source33(spike_out_source[33]),        .spike_out_source34(spike_out_source[34]),        .spike_out_source35(spike_out_source[35]),        .spike_out_source36(spike_out_source[36]),        .spike_out_source37(spike_out_source[37]),        .spike_out_source38(spike_out_source[38]),        .spike_out_source39(spike_out_source[39]),        .spike_out_source40(spike_out_source[40]),        .spike_out_source41(spike_out_source[41]),        .spike_out_source42(spike_out_source[42]),        .spike_out_source43(spike_out_source[43]),        .spike_out_source44(spike_out_source[44]),        .spike_out_source45(spike_out_source[45]),        .spike_out_source46(spike_out_source[46]),        .spike_out_source47(spike_out_source[47]),        .spike_out_source48(spike_out_source[48]),        .spike_out_source49(spike_out_source[49]),        .spike_out_source50(spike_out_source[50]),        .spike_out_source51(spike_out_source[51]),        .spike_out_source52(spike_out_source[52]),        .spike_out_source53(spike_out_source[53]),        .spike_out_source54(spike_out_source[54]),        .spike_out_source55(spike_out_source[55]),        .spike_out_source56(spike_out_source[56]),        .spike_out_source57(spike_out_source[57]),        .spike_out_source58(spike_out_source[58]),        .spike_out_source59(spike_out_source[59]),        .spike_out_source60(spike_out_source[60]),        .spike_out_source61(spike_out_source[61]),        .spike_out_source62(spike_out_source[62]),        .spike_out_source63(spike_out_source[63]),        .spike_out_source64(spike_out_source[64]),        .spike_out_source65(spike_out_source[65]),        .spike_out_source66(spike_out_source[66]),        .spike_out_source67(spike_out_source[67]),        .spike_out_source68(spike_out_source[68]),        .spike_out_source69(spike_out_source[69]),        .spike_out_source70(spike_out_source[70]),        .spike_out_source71(spike_out_source[71]),        .spike_out_source72(spike_out_source[72]),        .spike_out_source73(spike_out_source[73]),        .spike_out_source74(spike_out_source[74]),        .spike_out_source75(spike_out_source[75]),        .spike_out_source76(spike_out_source[76]),        .spike_out_source77(spike_out_source[77]),        .spike_out_source78(spike_out_source[78]),        .spike_out_source79(spike_out_source[79]),        .spike_out_source80(spike_out_source[80]),        .spike_out_source81(spike_out_source[81]),        .spike_out_source82(spike_out_source[82]),        .spike_out_source83(spike_out_source[83]),        .spike_out_source84(spike_out_source[84]),        .spike_out_source85(spike_out_source[85]),        .spike_out_source86(spike_out_source[86]),        .spike_out_source87(spike_out_source[87]),        .spike_out_source88(spike_out_source[88]),        .spike_out_source89(spike_out_source[89]),        .spike_out_source90(spike_out_source[90]),        .spike_out_source91(spike_out_source[91]),        .spike_out_source92(spike_out_source[92]),        .spike_out_source93(spike_out_source[93]),        .spike_out_source94(spike_out_source[94]),        .spike_out_source95(spike_out_source[95]),        .spike_out_source96(spike_out_source[96]),        .spike_out_source97(spike_out_source[97]),        .spike_out_source98(spike_out_source[98]),        .spike_out_source99(spike_out_source[99]),        .spike_out_source100(spike_out_source[100]),
        .spike_out_source101(spike_out_source[101]),        .spike_out_source102(spike_out_source[102]),        .spike_out_source103(spike_out_source[103]),        .spike_out_source104(spike_out_source[104]),        .spike_out_source105(spike_out_source[105]),        .spike_out_source106(spike_out_source[106]),        .spike_out_source107(spike_out_source[107]),        .spike_out_source108(spike_out_source[108]),        .spike_out_source109(spike_out_source[109]),        .spike_out_source110(spike_out_source[110]),        .spike_out_source111(spike_out_source[111]),        .spike_out_source112(spike_out_source[112]),        .spike_out_source113(spike_out_source[113]),        .spike_out_source114(spike_out_source[114]),        .spike_out_source115(spike_out_source[115]),        .spike_out_source116(spike_out_source[116]),        .spike_out_source117(spike_out_source[117]),        .spike_out_source118(spike_out_source[118]),        .spike_out_source119(spike_out_source[119]),        .spike_out_source120(spike_out_source[120]),        .spike_out_source121(spike_out_source[121]),        .spike_out_source122(spike_out_source[122]),        .spike_out_source123(spike_out_source[123]),        .spike_out_source124(spike_out_source[124]),        .spike_out_source125(spike_out_source[125]),        .spike_out_source126(spike_out_source[126]),        .spike_out_source127(spike_out_source[127]),        .spike_out_source128(spike_out_source[128]),        .spike_out_source129(spike_out_source[129]),        .spike_out_source130(spike_out_source[130]),        .spike_out_source131(spike_out_source[131]),        .spike_out_source132(spike_out_source[132]),        .spike_out_source133(spike_out_source[133]),        .spike_out_source134(spike_out_source[134]),        .spike_out_source135(spike_out_source[135]),        .spike_out_source136(spike_out_source[136]),        .spike_out_source137(spike_out_source[137]),        .spike_out_source138(spike_out_source[138]),        .spike_out_source139(spike_out_source[139]),        .spike_out_source140(spike_out_source[140]),        .spike_out_source141(spike_out_source[141]),        .spike_out_source142(spike_out_source[142]),        .spike_out_source143(spike_out_source[143]),        .spike_out_source144(spike_out_source[144]),        .spike_out_source145(spike_out_source[145]),        .spike_out_source146(spike_out_source[146]),        .spike_out_source147(spike_out_source[147]),        .spike_out_source148(spike_out_source[148]),        .spike_out_source149(spike_out_source[149]),        .spike_out_source150(spike_out_source[150]),        .spike_out_source151(spike_out_source[151]),        .spike_out_source152(spike_out_source[152]),        .spike_out_source153(spike_out_source[153]),        .spike_out_source154(spike_out_source[154]),        .spike_out_source155(spike_out_source[155]),        .spike_out_source156(spike_out_source[156]),        .spike_out_source157(spike_out_source[157]),        .spike_out_source158(spike_out_source[158]),        .spike_out_source159(spike_out_source[159]),        .spike_out_source160(spike_out_source[160]),        .spike_out_source161(spike_out_source[161]),        .spike_out_source162(spike_out_source[162]),        .spike_out_source163(spike_out_source[163]),        .spike_out_source164(spike_out_source[164]),        .spike_out_source165(spike_out_source[165]),        .spike_out_source166(spike_out_source[166]),        .spike_out_source167(spike_out_source[167]),        .spike_out_source168(spike_out_source[168]),        .spike_out_source169(spike_out_source[169]),        .spike_out_source170(spike_out_source[170]),        .spike_out_source171(spike_out_source[171]),        .spike_out_source172(spike_out_source[172]),        .spike_out_source173(spike_out_source[173]),        .spike_out_source174(spike_out_source[174]),        .spike_out_source175(spike_out_source[175]),        .spike_out_source176(spike_out_source[176]),        .spike_out_source177(spike_out_source[177]),        .spike_out_source178(spike_out_source[178]),        .spike_out_source179(spike_out_source[179]),        .spike_out_source180(spike_out_source[180]),        .spike_out_source181(spike_out_source[181]),        .spike_out_source182(spike_out_source[182]),        .spike_out_source183(spike_out_source[183]),        .spike_out_source184(spike_out_source[184]),        .spike_out_source185(spike_out_source[185]),        .spike_out_source186(spike_out_source[186]),        .spike_out_source187(spike_out_source[187]),        .spike_out_source188(spike_out_source[188]),        .spike_out_source189(spike_out_source[189]),        .spike_out_source190(spike_out_source[190]),        .spike_out_source191(spike_out_source[191]),        .spike_out_source192(spike_out_source[192]),        .spike_out_source193(spike_out_source[193]),        .spike_out_source194(spike_out_source[194]),        .spike_out_source195(spike_out_source[195]),        .spike_out_source196(spike_out_source[196]),        .spike_out_source197(spike_out_source[197]),        .spike_out_source198(spike_out_source[198]),        .spike_out_source199(spike_out_source[199]),        .spike_out_source200(spike_out_source[200]),
        .spike_out_source201(spike_out_source[201]),        .spike_out_source202(spike_out_source[202]),        .spike_out_source203(spike_out_source[203]),        .spike_out_source204(spike_out_source[204]),        .spike_out_source205(spike_out_source[205]),        .spike_out_source206(spike_out_source[206]),        .spike_out_source207(spike_out_source[207]),        .spike_out_source208(spike_out_source[208]),        .spike_out_source209(spike_out_source[209]),        .spike_out_source210(spike_out_source[210]),        .spike_out_source211(spike_out_source[211]),        .spike_out_source212(spike_out_source[212]),        .spike_out_source213(spike_out_source[213]),        .spike_out_source214(spike_out_source[214]),        .spike_out_source215(spike_out_source[215]),        .spike_out_source216(spike_out_source[216]),        .spike_out_source217(spike_out_source[217]),        .spike_out_source218(spike_out_source[218]),        .spike_out_source219(spike_out_source[219]),        .spike_out_source220(spike_out_source[220]),        .spike_out_source221(spike_out_source[221]),        .spike_out_source222(spike_out_source[222]),        .spike_out_source223(spike_out_source[223]),        .spike_out_source224(spike_out_source[224]),        .spike_out_source225(spike_out_source[225]),        .spike_out_source226(spike_out_source[226]),        .spike_out_source227(spike_out_source[227]),        .spike_out_source228(spike_out_source[228]),        .spike_out_source229(spike_out_source[229]),        .spike_out_source230(spike_out_source[230]),        .spike_out_source231(spike_out_source[231]),        .spike_out_source232(spike_out_source[232]),        .spike_out_source233(spike_out_source[233]),        .spike_out_source234(spike_out_source[234]),        .spike_out_source235(spike_out_source[235]),        .spike_out_source236(spike_out_source[236]),        .spike_out_source237(spike_out_source[237]),        .spike_out_source238(spike_out_source[238]),        .spike_out_source239(spike_out_source[239]),        .spike_out_source240(spike_out_source[240]),        .spike_out_source241(spike_out_source[241]),        .spike_out_source242(spike_out_source[242]),        .spike_out_source243(spike_out_source[243]),        .spike_out_source244(spike_out_source[244]),        .spike_out_source245(spike_out_source[245]),        .spike_out_source246(spike_out_source[246]),        .spike_out_source247(spike_out_source[247]),        .spike_out_source248(spike_out_source[248]),        .spike_out_source249(spike_out_source[249]),        .spike_out_source250(spike_out_source[250]),        .spike_out_source251(spike_out_source[251]),        .spike_out_source252(spike_out_source[252]),        .spike_out_source253(spike_out_source[253]),        .spike_out_source254(spike_out_source[254]),        .spike_out_source255(spike_out_source[255]),        .spike_out_source256(spike_out_source[256]),        .spike_out_source257(spike_out_source[257]),        .spike_out_source258(spike_out_source[258]),        .spike_out_source259(spike_out_source[259]),        .spike_out_source260(spike_out_source[260]),        .spike_out_source261(spike_out_source[261]),        .spike_out_source262(spike_out_source[262]),        .spike_out_source263(spike_out_source[263]),        .spike_out_source264(spike_out_source[264]),        .spike_out_source265(spike_out_source[265]),        .spike_out_source266(spike_out_source[266]),        .spike_out_source267(spike_out_source[267]),        .spike_out_source268(spike_out_source[268]),        .spike_out_source269(spike_out_source[269]),        .spike_out_source270(spike_out_source[270]),        .spike_out_source271(spike_out_source[271]),        .spike_out_source272(spike_out_source[272]),        .spike_out_source273(spike_out_source[273]),        .spike_out_source274(spike_out_source[274]),        .spike_out_source275(spike_out_source[275]),        .spike_out_source276(spike_out_source[276]),        .spike_out_source277(spike_out_source[277]),        .spike_out_source278(spike_out_source[278]),        .spike_out_source279(spike_out_source[279]),        .spike_out_source280(spike_out_source[280]),        .spike_out_source281(spike_out_source[281]),        .spike_out_source282(spike_out_source[282]),        .spike_out_source283(spike_out_source[283]),        .spike_out_source284(spike_out_source[284]),        .spike_out_source285(spike_out_source[285]),        .spike_out_source286(spike_out_source[286]),        .spike_out_source287(spike_out_source[287]),        .spike_out_source288(spike_out_source[288]),        .spike_out_source289(spike_out_source[289]),        .spike_out_source290(spike_out_source[290]),        .spike_out_source291(spike_out_source[291]),        .spike_out_source292(spike_out_source[292]),        .spike_out_source293(spike_out_source[293]),        .spike_out_source294(spike_out_source[294]),        .spike_out_source295(spike_out_source[295]),        .spike_out_source296(spike_out_source[296]),        .spike_out_source297(spike_out_source[297]),        .spike_out_source298(spike_out_source[298]),        .spike_out_source299(spike_out_source[299]),        .spike_out_source300(spike_out_source[300]),
        .spike_out_source301(spike_out_source[301]),        .spike_out_source302(spike_out_source[302]),        .spike_out_source303(spike_out_source[303]),        .spike_out_source304(spike_out_source[304]),        .spike_out_source305(spike_out_source[305]),        .spike_out_source306(spike_out_source[306]),        .spike_out_source307(spike_out_source[307]),        .spike_out_source308(spike_out_source[308]),        .spike_out_source309(spike_out_source[309]),        .spike_out_source310(spike_out_source[310]),        .spike_out_source311(spike_out_source[311]),        .spike_out_source312(spike_out_source[312]),        .spike_out_source313(spike_out_source[313]),        .spike_out_source314(spike_out_source[314]),        .spike_out_source315(spike_out_source[315]),        .spike_out_source316(spike_out_source[316]),        .spike_out_source317(spike_out_source[317]),        .spike_out_source318(spike_out_source[318]),        .spike_out_source319(spike_out_source[319]),        .spike_out_source320(spike_out_source[320]),        .spike_out_source321(spike_out_source[321]),        .spike_out_source322(spike_out_source[322]),        .spike_out_source323(spike_out_source[323]),        .spike_out_source324(spike_out_source[324]),        .spike_out_source325(spike_out_source[325]),        .spike_out_source326(spike_out_source[326]),        .spike_out_source327(spike_out_source[327]),        .spike_out_source328(spike_out_source[328]),        .spike_out_source329(spike_out_source[329]),        .spike_out_source330(spike_out_source[330]),        .spike_out_source331(spike_out_source[331]),        .spike_out_source332(spike_out_source[332]),        .spike_out_source333(spike_out_source[333]),        .spike_out_source334(spike_out_source[334]),        .spike_out_source335(spike_out_source[335]),        .spike_out_source336(spike_out_source[336]),        .spike_out_source337(spike_out_source[337]),        .spike_out_source338(spike_out_source[338]),        .spike_out_source339(spike_out_source[339]),        .spike_out_source340(spike_out_source[340]),        .spike_out_source341(spike_out_source[341]),        .spike_out_source342(spike_out_source[342]),        .spike_out_source343(spike_out_source[343]),        .spike_out_source344(spike_out_source[344]),        .spike_out_source345(spike_out_source[345]),        .spike_out_source346(spike_out_source[346]),        .spike_out_source347(spike_out_source[347]),        .spike_out_source348(spike_out_source[348]),        .spike_out_source349(spike_out_source[349]),        .spike_out_source350(spike_out_source[350]),        .spike_out_source351(spike_out_source[351]),        .spike_out_source352(spike_out_source[352]),        .spike_out_source353(spike_out_source[353]),        .spike_out_source354(spike_out_source[354]),        .spike_out_source355(spike_out_source[355]),        .spike_out_source356(spike_out_source[356]),        .spike_out_source357(spike_out_source[357]),        .spike_out_source358(spike_out_source[358]),        .spike_out_source359(spike_out_source[359]),        .spike_out_source360(spike_out_source[360]),        .spike_out_source361(spike_out_source[361]),        .spike_out_source362(spike_out_source[362]),        .spike_out_source363(spike_out_source[363]),        .spike_out_source364(spike_out_source[364]),        .spike_out_source365(spike_out_source[365]),        .spike_out_source366(spike_out_source[366]),        .spike_out_source367(spike_out_source[367]),        .spike_out_source368(spike_out_source[368]),        .spike_out_source369(spike_out_source[369]),        .spike_out_source370(spike_out_source[370]),        .spike_out_source371(spike_out_source[371]),        .spike_out_source372(spike_out_source[372]),        .spike_out_source373(spike_out_source[373]),        .spike_out_source374(spike_out_source[374]),        .spike_out_source375(spike_out_source[375]),        .spike_out_source376(spike_out_source[376]),        .spike_out_source377(spike_out_source[377]),        .spike_out_source378(spike_out_source[378]),        .spike_out_source379(spike_out_source[379]),        .spike_out_source380(spike_out_source[380]),        .spike_out_source381(spike_out_source[381]),        .spike_out_source382(spike_out_source[382]),        .spike_out_source383(spike_out_source[383]),        .spike_out_source384(spike_out_source[384]),        .spike_out_source385(spike_out_source[385]),        .spike_out_source386(spike_out_source[386]),        .spike_out_source387(spike_out_source[387]),        .spike_out_source388(spike_out_source[388]),        .spike_out_source389(spike_out_source[389]),        .spike_out_source390(spike_out_source[390]),        .spike_out_source391(spike_out_source[391]),        .spike_out_source392(spike_out_source[392]),        .spike_out_source393(spike_out_source[393]),        .spike_out_source394(spike_out_source[394]),        .spike_out_source395(spike_out_source[395]),        .spike_out_source396(spike_out_source[396]),        .spike_out_source397(spike_out_source[397]),        .spike_out_source398(spike_out_source[398]),        .spike_out_source399(spike_out_source[399]),        .spike_out_source400(spike_out_source[400]),
        .spike_out_source401(spike_out_source[401]),        .spike_out_source402(spike_out_source[402]),        .spike_out_source403(spike_out_source[403]),        .spike_out_source404(spike_out_source[404]),        .spike_out_source405(spike_out_source[405]),        .spike_out_source406(spike_out_source[406]),        .spike_out_source407(spike_out_source[407]),        .spike_out_source408(spike_out_source[408]),        .spike_out_source409(spike_out_source[409]),        .spike_out_source410(spike_out_source[410]),        .spike_out_source411(spike_out_source[411]),        .spike_out_source412(spike_out_source[412]),        .spike_out_source413(spike_out_source[413]),        .spike_out_source414(spike_out_source[414]),        .spike_out_source415(spike_out_source[415]),        .spike_out_source416(spike_out_source[416]),        .spike_out_source417(spike_out_source[417]),        .spike_out_source418(spike_out_source[418]),        .spike_out_source419(spike_out_source[419]),        .spike_out_source420(spike_out_source[420]),        .spike_out_source421(spike_out_source[421]),        .spike_out_source422(spike_out_source[422]),        .spike_out_source423(spike_out_source[423]),        .spike_out_source424(spike_out_source[424]),        .spike_out_source425(spike_out_source[425]),        .spike_out_source426(spike_out_source[426]),        .spike_out_source427(spike_out_source[427]),        .spike_out_source428(spike_out_source[428]),        .spike_out_source429(spike_out_source[429]),        .spike_out_source430(spike_out_source[430]),        .spike_out_source431(spike_out_source[431]),        .spike_out_source432(spike_out_source[432]),        .spike_out_source433(spike_out_source[433]),        .spike_out_source434(spike_out_source[434]),        .spike_out_source435(spike_out_source[435]),        .spike_out_source436(spike_out_source[436]),        .spike_out_source437(spike_out_source[437]),        .spike_out_source438(spike_out_source[438]),        .spike_out_source439(spike_out_source[439]),        .spike_out_source440(spike_out_source[440]),        .spike_out_source441(spike_out_source[441]),        .spike_out_source442(spike_out_source[442]),        .spike_out_source443(spike_out_source[443]),        .spike_out_source444(spike_out_source[444]),        .spike_out_source445(spike_out_source[445]),        .spike_out_source446(spike_out_source[446]),        .spike_out_source447(spike_out_source[447]),        .spike_out_source448(spike_out_source[448]),        .spike_out_source449(spike_out_source[449]),        .spike_out_source450(spike_out_source[450]),        .spike_out_source451(spike_out_source[451]),        .spike_out_source452(spike_out_source[452]),        .spike_out_source453(spike_out_source[453]),        .spike_out_source454(spike_out_source[454]),        .spike_out_source455(spike_out_source[455]),        .spike_out_source456(spike_out_source[456]),        .spike_out_source457(spike_out_source[457]),        .spike_out_source458(spike_out_source[458]),        .spike_out_source459(spike_out_source[459]),        .spike_out_source460(spike_out_source[460]),        .spike_out_source461(spike_out_source[461]),        .spike_out_source462(spike_out_source[462]),        .spike_out_source463(spike_out_source[463]),        .spike_out_source464(spike_out_source[464]),        .spike_out_source465(spike_out_source[465]),        .spike_out_source466(spike_out_source[466]),        .spike_out_source467(spike_out_source[467]),        .spike_out_source468(spike_out_source[468]),        .spike_out_source469(spike_out_source[469]),        .spike_out_source470(spike_out_source[470]),        .spike_out_source471(spike_out_source[471]),        .spike_out_source472(spike_out_source[472]),        .spike_out_source473(spike_out_source[473]),        .spike_out_source474(spike_out_source[474]),        .spike_out_source475(spike_out_source[475]),        .spike_out_source476(spike_out_source[476]),        .spike_out_source477(spike_out_source[477]),        .spike_out_source478(spike_out_source[478]),        .spike_out_source479(spike_out_source[479]),        .spike_out_source480(spike_out_source[480]),        .spike_out_source481(spike_out_source[481]),        .spike_out_source482(spike_out_source[482]),        .spike_out_source483(spike_out_source[483]),        .spike_out_source484(spike_out_source[484]),        .spike_out_source485(spike_out_source[485]),        .spike_out_source486(spike_out_source[486]),        .spike_out_source487(spike_out_source[487]),        .spike_out_source488(spike_out_source[488]),        .spike_out_source489(spike_out_source[489]),        .spike_out_source490(spike_out_source[490]),        .spike_out_source491(spike_out_source[491]),        .spike_out_source492(spike_out_source[492]),        .spike_out_source493(spike_out_source[493]),        .spike_out_source494(spike_out_source[494]),        .spike_out_source495(spike_out_source[495]),        .spike_out_source496(spike_out_source[496]),        .spike_out_source497(spike_out_source[497]),        .spike_out_source498(spike_out_source[498]),        .spike_out_source499(spike_out_source[499]),        .spike_out_source500(spike_out_source[500]),
        .spike_out_source501(spike_out_source[501]),        .spike_out_source502(spike_out_source[502]),        .spike_out_source503(spike_out_source[503]),        .spike_out_source504(spike_out_source[504]),        .spike_out_source505(spike_out_source[505]),        .spike_out_source506(spike_out_source[506]),        .spike_out_source507(spike_out_source[507]),        .spike_out_source508(spike_out_source[508]),        .spike_out_source509(spike_out_source[509]),        .spike_out_source510(spike_out_source[510]),        .spike_out_source511(spike_out_source[511]),        .spike_out_source512(spike_out_source[512]),        .spike_out_source513(spike_out_source[513]),        .spike_out_source514(spike_out_source[514]),        .spike_out_source515(spike_out_source[515]),        .spike_out_source516(spike_out_source[516]),        .spike_out_source517(spike_out_source[517]),        .spike_out_source518(spike_out_source[518]),        .spike_out_source519(spike_out_source[519]),        .spike_out_source520(spike_out_source[520]),        .spike_out_source521(spike_out_source[521]),        .spike_out_source522(spike_out_source[522]),        .spike_out_source523(spike_out_source[523]),        .spike_out_source524(spike_out_source[524]),        .spike_out_source525(spike_out_source[525]),        .spike_out_source526(spike_out_source[526]),        .spike_out_source527(spike_out_source[527]),        .spike_out_source528(spike_out_source[528]),        .spike_out_source529(spike_out_source[529]),        .spike_out_source530(spike_out_source[530]),        .spike_out_source531(spike_out_source[531]),        .spike_out_source532(spike_out_source[532]),        .spike_out_source533(spike_out_source[533]),        .spike_out_source534(spike_out_source[534]),        .spike_out_source535(spike_out_source[535]),        .spike_out_source536(spike_out_source[536]),        .spike_out_source537(spike_out_source[537]),        .spike_out_source538(spike_out_source[538]),        .spike_out_source539(spike_out_source[539]),        .spike_out_source540(spike_out_source[540]),        .spike_out_source541(spike_out_source[541]),        .spike_out_source542(spike_out_source[542]),        .spike_out_source543(spike_out_source[543]),        .spike_out_source544(spike_out_source[544]),        .spike_out_source545(spike_out_source[545]),        .spike_out_source546(spike_out_source[546]),        .spike_out_source547(spike_out_source[547]),        .spike_out_source548(spike_out_source[548]),        .spike_out_source549(spike_out_source[549]),        .spike_out_source550(spike_out_source[550]),        .spike_out_source551(spike_out_source[551]),        .spike_out_source552(spike_out_source[552]),        .spike_out_source553(spike_out_source[553]),        .spike_out_source554(spike_out_source[554]),        .spike_out_source555(spike_out_source[555]),        .spike_out_source556(spike_out_source[556]),        .spike_out_source557(spike_out_source[557]),        .spike_out_source558(spike_out_source[558]),        .spike_out_source559(spike_out_source[559]),        .spike_out_source560(spike_out_source[560]),        .spike_out_source561(spike_out_source[561]),        .spike_out_source562(spike_out_source[562]),        .spike_out_source563(spike_out_source[563]),        .spike_out_source564(spike_out_source[564]),        .spike_out_source565(spike_out_source[565]),        .spike_out_source566(spike_out_source[566]),        .spike_out_source567(spike_out_source[567]),        .spike_out_source568(spike_out_source[568]),        .spike_out_source569(spike_out_source[569]),        .spike_out_source570(spike_out_source[570]),        .spike_out_source571(spike_out_source[571]),        .spike_out_source572(spike_out_source[572]),        .spike_out_source573(spike_out_source[573]),        .spike_out_source574(spike_out_source[574]),        .spike_out_source575(spike_out_source[575]),        .spike_out_source576(spike_out_source[576]),        .spike_out_source577(spike_out_source[577]),        .spike_out_source578(spike_out_source[578]),        .spike_out_source579(spike_out_source[579]),        .spike_out_source580(spike_out_source[580]),        .spike_out_source581(spike_out_source[581]),        .spike_out_source582(spike_out_source[582]),        .spike_out_source583(spike_out_source[583]),        .spike_out_source584(spike_out_source[584]),        .spike_out_source585(spike_out_source[585]),        .spike_out_source586(spike_out_source[586]),        .spike_out_source587(spike_out_source[587]),        .spike_out_source588(spike_out_source[588]),        .spike_out_source589(spike_out_source[589]),        .spike_out_source590(spike_out_source[590]),        .spike_out_source591(spike_out_source[591]),        .spike_out_source592(spike_out_source[592]),        .spike_out_source593(spike_out_source[593]),        .spike_out_source594(spike_out_source[594]),        .spike_out_source595(spike_out_source[595]),        .spike_out_source596(spike_out_source[596]),        .spike_out_source597(spike_out_source[597]),        .spike_out_source598(spike_out_source[598]),        .spike_out_source599(spike_out_source[599]),        .spike_out_source600(spike_out_source[600]),
        .spike_out_source601(spike_out_source[601]),        .spike_out_source602(spike_out_source[602]),        .spike_out_source603(spike_out_source[603]),        .spike_out_source604(spike_out_source[604]),        .spike_out_source605(spike_out_source[605]),        .spike_out_source606(spike_out_source[606]),        .spike_out_source607(spike_out_source[607]),        .spike_out_source608(spike_out_source[608]),        .spike_out_source609(spike_out_source[609]),        .spike_out_source610(spike_out_source[610]),        .spike_out_source611(spike_out_source[611]),        .spike_out_source612(spike_out_source[612]),        .spike_out_source613(spike_out_source[613]),        .spike_out_source614(spike_out_source[614]),        .spike_out_source615(spike_out_source[615]),        .spike_out_source616(spike_out_source[616]),        .spike_out_source617(spike_out_source[617]),        .spike_out_source618(spike_out_source[618]),        .spike_out_source619(spike_out_source[619]),        .spike_out_source620(spike_out_source[620]),        .spike_out_source621(spike_out_source[621]),        .spike_out_source622(spike_out_source[622]),        .spike_out_source623(spike_out_source[623]),        .spike_out_source624(spike_out_source[624]),        .spike_out_source625(spike_out_source[625]),        .spike_out_source626(spike_out_source[626]),        .spike_out_source627(spike_out_source[627]),        .spike_out_source628(spike_out_source[628]),        .spike_out_source629(spike_out_source[629]),        .spike_out_source630(spike_out_source[630]),        .spike_out_source631(spike_out_source[631]),        .spike_out_source632(spike_out_source[632]),        .spike_out_source633(spike_out_source[633]),        .spike_out_source634(spike_out_source[634]),        .spike_out_source635(spike_out_source[635]),        .spike_out_source636(spike_out_source[636]),        .spike_out_source637(spike_out_source[637]),        .spike_out_source638(spike_out_source[638]),        .spike_out_source639(spike_out_source[639]),        .spike_out_source640(spike_out_source[640]),        .spike_out_source641(spike_out_source[641]),        .spike_out_source642(spike_out_source[642]),        .spike_out_source643(spike_out_source[643]),        .spike_out_source644(spike_out_source[644]),        .spike_out_source645(spike_out_source[645]),        .spike_out_source646(spike_out_source[646]),        .spike_out_source647(spike_out_source[647]),        .spike_out_source648(spike_out_source[648]),        .spike_out_source649(spike_out_source[649]),        .spike_out_source650(spike_out_source[650]),        .spike_out_source651(spike_out_source[651]),        .spike_out_source652(spike_out_source[652]),        .spike_out_source653(spike_out_source[653]),        .spike_out_source654(spike_out_source[654]),        .spike_out_source655(spike_out_source[655]),        .spike_out_source656(spike_out_source[656]),        .spike_out_source657(spike_out_source[657]),        .spike_out_source658(spike_out_source[658]),        .spike_out_source659(spike_out_source[659]),        .spike_out_source660(spike_out_source[660]),        .spike_out_source661(spike_out_source[661]),        .spike_out_source662(spike_out_source[662]),        .spike_out_source663(spike_out_source[663]),        .spike_out_source664(spike_out_source[664]),        .spike_out_source665(spike_out_source[665]),        .spike_out_source666(spike_out_source[666]),        .spike_out_source667(spike_out_source[667]),        .spike_out_source668(spike_out_source[668]),        .spike_out_source669(spike_out_source[669]),        .spike_out_source670(spike_out_source[670]),        .spike_out_source671(spike_out_source[671]),        .spike_out_source672(spike_out_source[672]),        .spike_out_source673(spike_out_source[673]),        .spike_out_source674(spike_out_source[674]),        .spike_out_source675(spike_out_source[675]),        .spike_out_source676(spike_out_source[676]),        .spike_out_source677(spike_out_source[677]),        .spike_out_source678(spike_out_source[678]),        .spike_out_source679(spike_out_source[679]),        .spike_out_source680(spike_out_source[680]),        .spike_out_source681(spike_out_source[681]),        .spike_out_source682(spike_out_source[682]),        .spike_out_source683(spike_out_source[683]),        .spike_out_source684(spike_out_source[684]),        .spike_out_source685(spike_out_source[685]),        .spike_out_source686(spike_out_source[686]),        .spike_out_source687(spike_out_source[687]),        .spike_out_source688(spike_out_source[688]),        .spike_out_source689(spike_out_source[689]),        .spike_out_source690(spike_out_source[690]),        .spike_out_source691(spike_out_source[691]),        .spike_out_source692(spike_out_source[692]),        .spike_out_source693(spike_out_source[693]),        .spike_out_source694(spike_out_source[694]),        .spike_out_source695(spike_out_source[695]),        .spike_out_source696(spike_out_source[696]),        .spike_out_source697(spike_out_source[697]),        .spike_out_source698(spike_out_source[698]),        .spike_out_source699(spike_out_source[699]),        .spike_out_source700(spike_out_source[700]),
        .spike_out_source701(spike_out_source[701]),        .spike_out_source702(spike_out_source[702]),        .spike_out_source703(spike_out_source[703]),        .spike_out_source704(spike_out_source[704]),        .spike_out_source705(spike_out_source[705]),        .spike_out_source706(spike_out_source[706]),        .spike_out_source707(spike_out_source[707]),        .spike_out_source708(spike_out_source[708]),        .spike_out_source709(spike_out_source[709]),        .spike_out_source710(spike_out_source[710]),        .spike_out_source711(spike_out_source[711]),        .spike_out_source712(spike_out_source[712]),        .spike_out_source713(spike_out_source[713]),        .spike_out_source714(spike_out_source[714]),        .spike_out_source715(spike_out_source[715]),        .spike_out_source716(spike_out_source[716]),        .spike_out_source717(spike_out_source[717]),        .spike_out_source718(spike_out_source[718]),        .spike_out_source719(spike_out_source[719]),        .spike_out_source720(spike_out_source[720]),        .spike_out_source721(spike_out_source[721]),        .spike_out_source722(spike_out_source[722]),        .spike_out_source723(spike_out_source[723]),        .spike_out_source724(spike_out_source[724]),        .spike_out_source725(spike_out_source[725]),        .spike_out_source726(spike_out_source[726]),        .spike_out_source727(spike_out_source[727]),        .spike_out_source728(spike_out_source[728]),        .spike_out_source729(spike_out_source[729]),        .spike_out_source730(spike_out_source[730]),        .spike_out_source731(spike_out_source[731]),        .spike_out_source732(spike_out_source[732]),        .spike_out_source733(spike_out_source[733]),        .spike_out_source734(spike_out_source[734]),        .spike_out_source735(spike_out_source[735]),        .spike_out_source736(spike_out_source[736]),        .spike_out_source737(spike_out_source[737]),        .spike_out_source738(spike_out_source[738]),        .spike_out_source739(spike_out_source[739]),        .spike_out_source740(spike_out_source[740]),        .spike_out_source741(spike_out_source[741]),        .spike_out_source742(spike_out_source[742]),        .spike_out_source743(spike_out_source[743]),        .spike_out_source744(spike_out_source[744]),        .spike_out_source745(spike_out_source[745]),        .spike_out_source746(spike_out_source[746]),        .spike_out_source747(spike_out_source[747]),        .spike_out_source748(spike_out_source[748]),        .spike_out_source749(spike_out_source[749]),        .spike_out_source750(spike_out_source[750]),        .spike_out_source751(spike_out_source[751]),        .spike_out_source752(spike_out_source[752]),        .spike_out_source753(spike_out_source[753]),        .spike_out_source754(spike_out_source[754]),        .spike_out_source755(spike_out_source[755]),        .spike_out_source756(spike_out_source[756]),        .spike_out_source757(spike_out_source[757]),        .spike_out_source758(spike_out_source[758]),        .spike_out_source759(spike_out_source[759]),        .spike_out_source760(spike_out_source[760]),        .spike_out_source761(spike_out_source[761]),        .spike_out_source762(spike_out_source[762]),        .spike_out_source763(spike_out_source[763]),        .spike_out_source764(spike_out_source[764]),        .spike_out_source765(spike_out_source[765]),        .spike_out_source766(spike_out_source[766]),        .spike_out_source767(spike_out_source[767]),        .spike_out_source768(spike_out_source[768]),        .spike_out_source769(spike_out_source[769]),        .spike_out_source770(spike_out_source[770]),        .spike_out_source771(spike_out_source[771]),        .spike_out_source772(spike_out_source[772]),        .spike_out_source773(spike_out_source[773]),        .spike_out_source774(spike_out_source[774]),        .spike_out_source775(spike_out_source[775]),        .spike_out_source776(spike_out_source[776]),        .spike_out_source777(spike_out_source[777]),        .spike_out_source778(spike_out_source[778]),        .spike_out_source779(spike_out_source[779]),        .spike_out_source780(spike_out_source[780]),        .spike_out_source781(spike_out_source[781]),        .spike_out_source782(spike_out_source[782]),        .spike_out_source783(spike_out_source[783]),        .spike_out_source784(spike_out_source[784]),        .spike_out_source785(spike_out_source[785]),        .spike_out_source786(spike_out_source[786]),        .spike_out_source787(spike_out_source[787]),        .spike_out_source788(spike_out_source[788]),        .spike_out_source789(spike_out_source[789]),        .spike_out_source790(spike_out_source[790]),        .spike_out_source791(spike_out_source[791]),        .spike_out_source792(spike_out_source[792]),        .spike_out_source793(spike_out_source[793]),        .spike_out_source794(spike_out_source[794]),        .spike_out_source795(spike_out_source[795]),        .spike_out_source796(spike_out_source[796]),        .spike_out_source797(spike_out_source[797]),        .spike_out_source798(spike_out_source[798]),        .spike_out_source799(spike_out_source[799]),        .spike_out_source800(spike_out_source[800]),
        .spike_out_source801(spike_out_source[801]),        .spike_out_source802(spike_out_source[802]),        .spike_out_source803(spike_out_source[803]),        .spike_out_source804(spike_out_source[804]),        .spike_out_source805(spike_out_source[805]),        .spike_out_source806(spike_out_source[806]),        .spike_out_source807(spike_out_source[807]),        .spike_out_source808(spike_out_source[808]),        .spike_out_source809(spike_out_source[809]),        .spike_out_source810(spike_out_source[810]),        .spike_out_source811(spike_out_source[811]),        .spike_out_source812(spike_out_source[812]),        .spike_out_source813(spike_out_source[813]),        .spike_out_source814(spike_out_source[814]),        .spike_out_source815(spike_out_source[815]),        .spike_out_source816(spike_out_source[816]),        .spike_out_source817(spike_out_source[817]),        .spike_out_source818(spike_out_source[818]),        .spike_out_source819(spike_out_source[819]),        .spike_out_source820(spike_out_source[820]),        .spike_out_source821(spike_out_source[821]),        .spike_out_source822(spike_out_source[822]),        .spike_out_source823(spike_out_source[823]),        .spike_out_source824(spike_out_source[824]),        .spike_out_source825(spike_out_source[825]),        .spike_out_source826(spike_out_source[826]),        .spike_out_source827(spike_out_source[827]),        .spike_out_source828(spike_out_source[828]),        .spike_out_source829(spike_out_source[829]),        .spike_out_source830(spike_out_source[830]),        .spike_out_source831(spike_out_source[831]),        .spike_out_source832(spike_out_source[832]),        .spike_out_source833(spike_out_source[833]),        .spike_out_source834(spike_out_source[834]),        .spike_out_source835(spike_out_source[835]),        .spike_out_source836(spike_out_source[836]),        .spike_out_source837(spike_out_source[837]),        .spike_out_source838(spike_out_source[838]),        .spike_out_source839(spike_out_source[839]),        .spike_out_source840(spike_out_source[840]),        .spike_out_source841(spike_out_source[841]),        .spike_out_source842(spike_out_source[842]),        .spike_out_source843(spike_out_source[843]),        .spike_out_source844(spike_out_source[844]),        .spike_out_source845(spike_out_source[845]),        .spike_out_source846(spike_out_source[846]),        .spike_out_source847(spike_out_source[847]),        .spike_out_source848(spike_out_source[848]),        .spike_out_source849(spike_out_source[849]),        .spike_out_source850(spike_out_source[850]),        .spike_out_source851(spike_out_source[851]),        .spike_out_source852(spike_out_source[852]),        .spike_out_source853(spike_out_source[853]),        .spike_out_source854(spike_out_source[854]),        .spike_out_source855(spike_out_source[855]),        .spike_out_source856(spike_out_source[856]),        .spike_out_source857(spike_out_source[857]),        .spike_out_source858(spike_out_source[858]),        .spike_out_source859(spike_out_source[859]),        .spike_out_source860(spike_out_source[860]),        .spike_out_source861(spike_out_source[861]),        .spike_out_source862(spike_out_source[862]),        .spike_out_source863(spike_out_source[863]),        .spike_out_source864(spike_out_source[864]),        .spike_out_source865(spike_out_source[865]),        .spike_out_source866(spike_out_source[866]),        .spike_out_source867(spike_out_source[867]),        .spike_out_source868(spike_out_source[868]),        .spike_out_source869(spike_out_source[869]),        .spike_out_source870(spike_out_source[870]),        .spike_out_source871(spike_out_source[871]),        .spike_out_source872(spike_out_source[872]),        .spike_out_source873(spike_out_source[873]),        .spike_out_source874(spike_out_source[874]),        .spike_out_source875(spike_out_source[875]),        .spike_out_source876(spike_out_source[876]),        .spike_out_source877(spike_out_source[877]),        .spike_out_source878(spike_out_source[878]),        .spike_out_source879(spike_out_source[879]),        .spike_out_source880(spike_out_source[880]),        .spike_out_source881(spike_out_source[881]),        .spike_out_source882(spike_out_source[882]),        .spike_out_source883(spike_out_source[883]),        .spike_out_source884(spike_out_source[884]),        .spike_out_source885(spike_out_source[885]),        .spike_out_source886(spike_out_source[886]),        .spike_out_source887(spike_out_source[887]),        .spike_out_source888(spike_out_source[888]),        .spike_out_source889(spike_out_source[889]),        .spike_out_source890(spike_out_source[890]),        .spike_out_source891(spike_out_source[891]),        .spike_out_source892(spike_out_source[892]),        .spike_out_source893(spike_out_source[893]),        .spike_out_source894(spike_out_source[894]),        .spike_out_source895(spike_out_source[895]),        .spike_out_source896(spike_out_source[896]),        .spike_out_source897(spike_out_source[897]),        .spike_out_source898(spike_out_source[898]),        .spike_out_source899(spike_out_source[899]),        .spike_out_source900(spike_out_source[900]),
        .spike_out_source901(spike_out_source[901]),        .spike_out_source902(spike_out_source[902]),        .spike_out_source903(spike_out_source[903]),        .spike_out_source904(spike_out_source[904]),        .spike_out_source905(spike_out_source[905]),        .spike_out_source906(spike_out_source[906]),        .spike_out_source907(spike_out_source[907]),        .spike_out_source908(spike_out_source[908]),        .spike_out_source909(spike_out_source[909]),        .spike_out_source910(spike_out_source[910]),        .spike_out_source911(spike_out_source[911]),        .spike_out_source912(spike_out_source[912]),        .spike_out_source913(spike_out_source[913]),        .spike_out_source914(spike_out_source[914]),        .spike_out_source915(spike_out_source[915]),        .spike_out_source916(spike_out_source[916]),        .spike_out_source917(spike_out_source[917]),        .spike_out_source918(spike_out_source[918]),        .spike_out_source919(spike_out_source[919]),        .spike_out_source920(spike_out_source[920]),        .spike_out_source921(spike_out_source[921]),        .spike_out_source922(spike_out_source[922]),        .spike_out_source923(spike_out_source[923]),        .spike_out_source924(spike_out_source[924]),        .spike_out_source925(spike_out_source[925]),        .spike_out_source926(spike_out_source[926]),        .spike_out_source927(spike_out_source[927]),        .spike_out_source928(spike_out_source[928]),        .spike_out_source929(spike_out_source[929]),        .spike_out_source930(spike_out_source[930]),        .spike_out_source931(spike_out_source[931]),        .spike_out_source932(spike_out_source[932]),        .spike_out_source933(spike_out_source[933]),        .spike_out_source934(spike_out_source[934]),        .spike_out_source935(spike_out_source[935]),        .spike_out_source936(spike_out_source[936]),        .spike_out_source937(spike_out_source[937]),        .spike_out_source938(spike_out_source[938]),        .spike_out_source939(spike_out_source[939]),        .spike_out_source940(spike_out_source[940]),        .spike_out_source941(spike_out_source[941]),        .spike_out_source942(spike_out_source[942]),        .spike_out_source943(spike_out_source[943]),        .spike_out_source944(spike_out_source[944]),        .spike_out_source945(spike_out_source[945]),        .spike_out_source946(spike_out_source[946]),        .spike_out_source947(spike_out_source[947]),        .spike_out_source948(spike_out_source[948]),        .spike_out_source949(spike_out_source[949]),        .spike_out_source950(spike_out_source[950]),        .spike_out_source951(spike_out_source[951]),        .spike_out_source952(spike_out_source[952]),        .spike_out_source953(spike_out_source[953]),        .spike_out_source954(spike_out_source[954]),        .spike_out_source955(spike_out_source[955]),        .spike_out_source956(spike_out_source[956]),        .spike_out_source957(spike_out_source[957]),        .spike_out_source958(spike_out_source[958]),        .spike_out_source959(spike_out_source[959]),        .spike_out_source960(spike_out_source[960]),        .spike_out_source961(spike_out_source[961]),        .spike_out_source962(spike_out_source[962]),        .spike_out_source963(spike_out_source[963]),        .spike_out_source964(spike_out_source[964]),        .spike_out_source965(spike_out_source[965]),        .spike_out_source966(spike_out_source[966]),        .spike_out_source967(spike_out_source[967]),        .spike_out_source968(spike_out_source[968]),        .spike_out_source969(spike_out_source[969]),        .spike_out_source970(spike_out_source[970]),        .spike_out_source971(spike_out_source[971]),        .spike_out_source972(spike_out_source[972]),        .spike_out_source973(spike_out_source[973]),        .spike_out_source974(spike_out_source[974]),        .spike_out_source975(spike_out_source[975]),        .spike_out_source976(spike_out_source[976]),        .spike_out_source977(spike_out_source[977]),        .spike_out_source978(spike_out_source[978]),        .spike_out_source979(spike_out_source[979]),        .spike_out_source980(spike_out_source[980]),        .spike_out_source981(spike_out_source[981]),        .spike_out_source982(spike_out_source[982]),        .spike_out_source983(spike_out_source[983]),        .spike_out_source984(spike_out_source[984]),        .spike_out_source985(spike_out_source[985]),        .spike_out_source986(spike_out_source[986]),        .spike_out_source987(spike_out_source[987]),        .spike_out_source988(spike_out_source[988]),        .spike_out_source989(spike_out_source[989]),        .spike_out_source990(spike_out_source[990]),        .spike_out_source991(spike_out_source[991]),        .spike_out_source992(spike_out_source[992]),        .spike_out_source993(spike_out_source[993]),        .spike_out_source994(spike_out_source[994]),        .spike_out_source995(spike_out_source[995]),        .spike_out_source996(spike_out_source[996]),        .spike_out_source997(spike_out_source[997]),        .spike_out_source998(spike_out_source[998]),        .spike_out_source999(spike_out_source[999]),        .spike_out_source1000(spike_out_source[1000]),
        .spike_out_source1001(spike_out_source[1001]),        .spike_out_source1002(spike_out_source[1002]),        .spike_out_source1003(spike_out_source[1003]),        .spike_out_source1004(spike_out_source[1004]),        .spike_out_source1005(spike_out_source[1005]),        .spike_out_source1006(spike_out_source[1006]),        .spike_out_source1007(spike_out_source[1007]),        .spike_out_source1008(spike_out_source[1008]),        .spike_out_source1009(spike_out_source[1009]),        .spike_out_source1010(spike_out_source[1010]),        .spike_out_source1011(spike_out_source[1011]),        .spike_out_source1012(spike_out_source[1012]),        .spike_out_source1013(spike_out_source[1013]),        .spike_out_source1014(spike_out_source[1014]),        .spike_out_source1015(spike_out_source[1015]),        .spike_out_source1016(spike_out_source[1016]),        .spike_out_source1017(spike_out_source[1017]),        .spike_out_source1018(spike_out_source[1018]),        .spike_out_source1019(spike_out_source[1019]),        .spike_out_source1020(spike_out_source[1020]),        .spike_out_source1021(spike_out_source[1021]),        .spike_out_source1022(spike_out_source[1022]),        .spike_out_source1023(spike_out_source[1023])
    );

    // Observe the timing on gtkwave
    initial
    begin
        $dumpfile("testbench.vcd");
        $dumpvars(0, testbench);
    end

    // // Print the outputs when ever the inputs change
    initial
    begin
        $monitor($time, "  Neuron_address: %b\n                     Membrane Potential: %b\n                     Decay Rate: %d\n                     After Potential Decay: %b\n                     Source_address: %b\n                     MAC result: %b\n                     Threshold: %b\n                     Output Potential: %b\n                     Spiked:%b", neuron_addresses[0], membrane_potential[0], decay_rate, results_potential_decay[0], source_addresses[0], results_mac[0],v_threshold[0],final_potential[0], spike[0]);
    end

    // Observe the timing on gtkwave
    initial begin
        $dumpfile("accelerator_wavedata.vcd");
        $dumpvars(0,testbench);
    end


    initial begin

        CLK = 1'b0;
        CLK_count = 0;
        clear = 1'b0;

        // for async fifo
        rst_n = 0;
        wr_en = 0;
        rd_en = 0;

        //decay rate for potential decay calculation
        decay_rate = 4'b0010;

        //type of SNN model run
        model = 2'b00;

        //neuron addresses
        neuron_addresses[0] = 12'd0;
        neuron_addresses[1] = 12'd1;    neuron_addresses[2] = 12'd2;    neuron_addresses[3] = 12'd3;    neuron_addresses[4] = 12'd4;    neuron_addresses[5] = 12'd5;    neuron_addresses[6] = 12'd6;    neuron_addresses[7] = 12'd7;    neuron_addresses[8] = 12'd8;    neuron_addresses[9] = 12'd9;


        //for network interface
        neuron_addresses_initialization = {        neuron_addresses[0], 
        neuron_addresses[1],         neuron_addresses[2],         neuron_addresses[3],         neuron_addresses[4],         neuron_addresses[5],         neuron_addresses[6],         neuron_addresses[7],         neuron_addresses[8],         neuron_addresses[9]};

        //CSR
        connection_pointer_initialization = {5'd0, 5'd3, 5'd5, 5'd8, 5'd10, 5'd12, 5'd14, 5'd15, 5'd17, 5'd18, 5'd19};

        downstream_connections_initialization = {12'b000000000011, 12'b000000000101, 12'b000000000111, 
        12'b000000000100, 12'b000000000110,
        12'b000000000100, 12'b000000000101, 12'b000000000110,
        12'b000000001000, 12'b000000001001,
        12'b000000001000, 12'b000000001001,
        12'b000000001000, 12'b000000001001,
        12'b000000001001,
        12'b000000001000, 12'b000000001001,
        12'b111111111011,
        12'b111111111100,
        132'd0};

        //initial membrane potential values
        membrane_potential[0] = 32'h41deb852;
        membrane_potential[1] = 32'h42806b85;
        membrane_potential[2] = 32'h40b75c29;
        membrane_potential[3] = 32'h4228b852;
        membrane_potential[4] = 32'h42aeb852;
        membrane_potential[5] = 32'h429deb85;
        membrane_potential[6] = 32'h4165eb85;
        membrane_potential[7] = 32'h4212147b;
        membrane_potential[8] = 32'h428e2e14;
        membrane_potential[9] = 32'h411a147b;

        //send source addresses array first
        source_addresses_arrays[0] = {12'b001111111000, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111};
        source_addresses_arrays[1] = {12'd3, 12'd4, 12'd5, 12'd6, 12'd7};
        source_addresses_arrays[2] = {12'd3, 12'd4, 12'd5, 12'd6, 12'd7};
        source_addresses_arrays[3] = {12'd0, 12'd4, 12'd5, 12'd6, 12'd7};
        source_addresses_arrays[4] = {12'd1, 12'd2, 12'd5, 12'd0, 12'd0};
        source_addresses_arrays[5] = {12'd0, 12'd4, 12'd5, 12'd6, 12'd7};
        source_addresses_arrays[6] = {12'd3, 12'd4, 12'd5, 12'd6, 12'd7};
        source_addresses_arrays[7] = {12'd3, 12'd4, 12'd5, 12'd6, 12'd7};
        source_addresses_arrays[8] = {12'd3, 12'd4, 12'd5, 12'd6, 12'd7};
        source_addresses_arrays[9] = {12'd3, 12'd4, 12'd5, 12'd6, 12'd7};

        //assign the weights
        weights_arrays[0] = {32'h4290b333, 32'h41975c29, 32'h42470a3d, 32'h0, 32'h42ae3852};
        weights_arrays[1] = {32'h4290b333, 32'h41975c29, 32'h42470a3d, 32'h0, 32'h42ae3852};
        weights_arrays[2] = {32'h4290b333, 32'h41975c29, 32'h42470a3d, 32'h0, 32'h42ae3852};
        weights_arrays[3] = {32'h4290b333, 32'h41975c29, 32'h42470a3d, 32'h0, 32'h42ae3852};
        weights_arrays[4] = {32'h423f47ae, 32'h4109999a, 32'h0, 32'h0, 32'h0};
        weights_arrays[5] = {32'h4290b333, 32'h41975c29, 32'h42470a3d, 32'h0, 32'h42ae3852};
        weights_arrays[6] = {32'h4290b333, 32'h41975c29, 32'h42470a3d, 32'h0, 32'h42ae3852};
        weights_arrays[7] = {32'h4290b333, 32'h41975c29, 32'h42470a3d, 32'h0, 32'h42ae3852};
        weights_arrays[8] = {32'h4290b333, 32'h41975c29, 32'h42470a3d, 32'h0, 32'h42ae3852};
        weights_arrays[9] = {32'h4290b333, 32'h41975c29, 32'h42470a3d, 32'h0, 32'h42ae3852};

        //threshold values
        v_threshold[0] = 32'h42200000;
        v_threshold[1] = 32'h4237851f;
        v_threshold[2] = 32'h4048f5c3;
        v_threshold[3] = 32'h42910000;
        v_threshold[4] = 32'h43480000;
        v_threshold[5] = 32'h426b28f6;
        v_threshold[6] = 32'h42200000;
        v_threshold[7] = 32'h43480000;
        v_threshold[8] = 32'h4215ae14;
        v_threshold[9] = 32'h4287c7ae;

        //Izikeivich Parameters
        a = 32'h4287c7ae;
        b = 32'h4287c7ae;
        c = 32'h4287c7ae;
        d = 32'h4287c7ae;
        u_initialize = 32'h4287c7ae;

        // #40
        // spike_out_source[0] = 12'b001111111000;
        // source_addresses[1] = 12'd3;

        #1 rst_n = 1;

        #300
        $finish;

    end

    //when packets arrive from the potential adder send the source address to the relevant mac unit 
    // always @(packet1) begin
    //     spike_origin = packet1[23:12];               // From where the spike came
    //     spike_destination = packet1[11:0];           // To where it should be sent 

    //     source_addresses[spike_destination] = spike_origin;      // Trigger the wire of the relevant accumulator
    // end

    // always @(packet1) begin 
    //     spike_origin = packet1[23:12];
    //     spike_destination = packet1[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet2) begin 
    //     spike_origin = packet2[23:12];
    //     spike_destination = packet2[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet3) begin 
    //     spike_origin = packet3[23:12];
    //     spike_destination = packet3[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet4) begin 
    //     spike_origin = packet4[23:12];
    //     spike_destination = packet4[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet5) begin 
    //     spike_origin = packet5[23:12];
    //     spike_destination = packet5[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet6) begin 
    //     spike_origin = packet6[23:12];
    //     spike_destination = packet6[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet7) begin 
    //     spike_origin = packet7[23:12];
    //     spike_destination = packet7[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet8) begin 
    //     spike_origin = packet8[23:12];
    //     spike_destination = packet8[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet9) begin 
    //     spike_origin = packet9[23:12];
    //     spike_destination = packet9[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet10) begin 
    //     spike_origin = packet10[23:12];
    //     spike_destination = packet10[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet11) begin 
    //     spike_origin = packet11[23:12];
    //     spike_destination = packet11[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet12) begin 
    //     spike_origin = packet12[23:12];
    //     spike_destination = packet12[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet13) begin 
    //     spike_origin = packet13[23:12];
    //     spike_destination = packet13[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet14) begin 
    //     spike_origin = packet14[23:12];
    //     spike_destination = packet14[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet15) begin 
    //     spike_origin = packet15[23:12];
    //     spike_destination = packet15[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet16) begin 
    //     spike_origin = packet16[23:12];
    //     spike_destination = packet16[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet17) begin 
    //     spike_origin = packet17[23:12];
    //     spike_destination = packet17[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet18) begin 
    //     spike_origin = packet18[23:12];
    //     spike_destination = packet18[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet19) begin 
    //     spike_origin = packet19[23:12];
    //     spike_destination = packet19[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet20) begin 
    //     spike_origin = packet20[23:12];
    //     spike_destination = packet20[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end
    // always @(packet21) begin 
    //     spike_origin = packet21[23:12];
    //     spike_destination = packet21[11:0];
    //     source_addresses[spike_destination] = spike_origin;
    // end

    //invert clock every 4 seconds
    always
        #4 CLK = ~CLK;

    //timestep is 4 clockcycles
    always @(posedge CLK) begin

        if(CLK_count==3) begin
            CLK_count=0;
            clear = 1'b1;
            wr_en = 0;
        end else begin
            CLK_count = CLK_count+1;
        end

        if(CLK_count == 0) begin
            wr_en = 1;
        end

        if(CLK_count==1) begin
            clear = 1'b0;
            // rd_en = 0;
        end
    end


endmodule
