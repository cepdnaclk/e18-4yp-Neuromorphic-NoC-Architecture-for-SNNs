module testbench_scaled;

    //Initialize downstream connections
        connection_pointer_initialization = {        12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd784,         12'd785,         12'd786,         12'd787,         12'd788,         12'd789,         12'd790,         12'd791,         12'd792,         12'd793,         12'd794,         12'd795,         12'd796,         12'd797,         12'd798,         12'd799,         12'd800,         12'd801,         12'd802,         12'd803,         12'd804,         12'd805,         12'd806,         12'd807,         12'd808,         12'd809,         12'd810,         12'd811,         12'd812,         12'd813,         12'd814,         12'd815,         12'd816,         12'd817,         12'd818,         12'd819,         12'd820,         12'd821,         12'd822,         12'd823,         12'd824,         12'd825,         12'd826,         12'd827,         12'd828,         12'd829,         12'd830,         12'd831,         12'd832,         12'd833,         12'd834,         12'd835,         12'd836,         12'd837,         12'd838,         12'd839,         12'd840,         12'd841,         12'd842,         12'd843,         12'd844,         12'd845,         12'd846,         12'd847,         12'd848,         12'd849,         12'd850,         12'd851,         12'd852,         12'd853,         12'd854,         12'd855,         12'd856,         12'd857,         12'd858,         12'd859,         12'd860,         12'd861,         12'd862,         12'd863,         12'd864,         12'd865,         12'd866,         12'd867,         12'd868,         12'd869,         12'd870,         12'd871,         12'd872,         12'd873,         12'd874,         12'd875,         12'd876,         12'd877,         12'd878,         12'd879,         12'd880,         12'd881,         12'd882,         12'd883,         12'd884,         12'd885,         12'd886,         12'd887,         12'd888,         12'd889,         12'd890,         12'd891,         12'd892,         12'd893,         12'd894,         12'd895,         12'd896,         12'd897,         12'd898,         12'd899,         12'd900,         12'd901,         12'd902,         12'd903,         12'd904,         12'd905,         12'd906,         12'd907,         12'd908,         12'd909,         12'd910,         12'd911,         12'd912,         12'd913,         12'd914,         12'd915,         12'd916,         12'd917,         12'd918,         12'd919,         12'd920,         12'd921,         12'd922,         12'd923,         12'd924,         12'd925,         12'd926,         12'd927,         12'd928,         12'd929,         12'd930,         12'd931,         12'd932,         12'd933,         12'd934,         12'd935,         12'd936,         12'd937,         12'd938,         12'd939,         12'd940,         12'd941,         12'd942,         12'd943,         12'd944,         12'd945,         12'd946,         12'd947,         12'd948,         12'd949,         12'd950,         12'd951,         12'd952,         12'd953,         12'd954,         12'd955,         12'd956,         12'd957,         12'd958,         12'd959,         12'd960,         12'd961,         12'd962,         12'd963,         12'd964,         12'd965,         12'd966,         12'd967,         12'd968,         12'd969,         12'd970,         12'd971,         12'd972,         12'd973,         12'd974,         12'd975,         12'd976,         12'd977,         12'd978,         12'd979,         12'd980,         12'd981,         12'd982,         12'd983,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993,         12'd984,         12'd985,         12'd986,         12'd987,         12'd988,         12'd989,         12'd990,         12'd991,         12'd992,         12'd993};





endmodule
